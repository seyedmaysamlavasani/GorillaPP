module RREncode(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_1(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_2(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateGenerator(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_rankCalc_req_ready,
    output mainOff_rankCalc_req_valid,
    output[63:0] mainOff_rankCalc_req_bits_damping,
    output[63:0] mainOff_rankCalc_req_bits_rank,
    output[31:0] mainOff_rankCalc_req_bits_fanoutDegree,
    output[9:0] mainOff_rankCalc_req_tag,
    output mainOff_rankCalc_rep_ready,
    input  mainOff_rankCalc_rep_valid,
    input [63:0] mainOff_rankCalc_rep_bits_out,
    input [9:0] mainOff_rankCalc_rep_tag);

  wire memPort_req_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[4:0] T10;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T11;
  reg[0:0] subStateTh_1;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T15;
  wire AllOffloadsValid_1;
  wire T16;
  wire T17;
  wire T18;
  reg[0:0] rankCalcPortHadValidRequest_1;
  wire T19;
  wire T20;
  wire T21;
  wire rankCalcPort_req_valid;
  wire T22;
  wire T23;
  wire T24;
  wire[7:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg[0:0] rankCalc_valid_received_1;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[9:0] T35;
  wire[9:0] rankCalcPort_rep_tag;
  wire rankCalcPort_rep_ready;
  wire[9:0] rankCalcPort_req_tag;
  wire[9:0] T36;
  wire rankCalcPort_rep_valid;
  wire T37;
  wire T38;
  wire[4:0] T39;
  wire T40;
  wire T41;
  reg[0:0] rankCalc_valid_received_0;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[9:0] T46;
  wire T47;
  wire T48;
  wire[4:0] T49;
  wire T50;
  wire T51;
  wire[4:0] T52;
  wire T53;
  wire T54;
  wire[4:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[9:0] T59;
  wire T60;
  wire T61;
  reg[0:0] memPortHadValidRequest_1;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[4:0] T66;
  wire T67;
  wire T68;
  wire[4:0] T69;
  wire T70;
  reg[0:0] mem_valid_received_1;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[9:0] T75;
  wire[9:0] memPort_rep_tag;
  wire memPort_rep_valid;
  wire T76;
  wire T77;
  wire[4:0] T78;
  wire T79;
  wire T80;
  wire[9:0] T81;
  wire T82;
  wire T83;
  wire AllOffloadsValid_0;
  wire T84;
  wire T85;
  wire T86;
  reg[0:0] rankCalcPortHadValidRequest_0;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[4:0] T91;
  wire T92;
  wire T93;
  wire[4:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire[9:0] T98;
  wire T99;
  wire T100;
  reg[0:0] memPortHadValidRequest_0;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  wire[4:0] T108;
  wire T109;
  reg[0:0] mem_valid_received_0;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire[9:0] T114;
  wire T115;
  wire T116;
  wire[4:0] T117;
  wire T118;
  wire T119;
  wire[9:0] T120;
  wire T121;
  reg[0:0] subStateTh_0;
  wire T122;
  wire T123;
  wire T124;
  wire[1:0] T125;
  wire T126;
  wire T127;
  reg[7:0] State_0;
  wire T128;
  wire T129;
  wire T130;
  wire[1:0] T131;
  wire[4:0] T132;
  wire T133;
  wire T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[7:0] T137;
  wire[7:0] T138;
  wire T139;
  reg[7:0] State_1;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire[7:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[7:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire[7:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[31:0] page_fanoutDegree;
  wire[31:0] T165;
  wire[127:0] memRep1_data;
  wire[127:0] T166;
  wire[127:0] memPortReplyValue;
  wire[127:0] T167;
  wire[127:0] T168;
  wire[127:0] T169;
  wire[127:0] T170;
  reg[127:0] memPortReplyStorage_1_data;
  wire T171;
  wire T172;
  wire[1:0] T173;
  wire[1024:0] T174;
  wire[127:0] T175;
  wire[127:0] memPort_rep_bits_data;
  wire T176;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  reg[0:0] outputReg_1_done;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  reg[0:0] inputReg_1_done;
  wire T199;
  wire T200;
  wire[1:0] T201;
  wire[4:0] T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  reg[0:0] inputReg_0_done;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  reg[0:0] outputReg_0_done;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  reg[31:0] outputReg_1_pageId;
  wire T218;
  wire[31:0] T219;
  wire[31:0] T220;
  wire[31:0] T221;
  wire[31:0] T222;
  wire[31:0] T223;
  reg[31:0] pageId_1;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire[31:0] T229;
  wire[31:0] T230;
  wire[31:0] T231;
  wire[31:0] T232;
  wire[31:0] T233;
  reg[31:0] inputReg_1_length;
  wire[31:0] T234;
  wire[31:0] T235;
  wire[31:0] T236;
  reg[31:0] inputReg_0_length;
  wire[31:0] T237;
  wire[31:0] T238;
  wire[31:0] T239;
  wire[31:0] T240;
  reg[31:0] inputReg_1_startPageId;
  wire[31:0] T241;
  wire[31:0] T242;
  wire[31:0] T243;
  reg[31:0] inputReg_0_startPageId;
  wire[31:0] T244;
  wire T245;
  wire T246;
  wire[31:0] T247;
  wire[31:0] T248;
  wire[31:0] T249;
  reg[31:0] fanoutDegree_1;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire[7:0] T257;
  wire T258;
  wire T259;
  wire T260;
  wire[31:0] T261;
  wire[31:0] T262;
  wire[31:0] T263;
  wire[31:0] T264;
  wire[31:0] T265;
  reg[31:0] fanoutDegree_0;
  wire T266;
  wire T267;
  wire T268;
  wire[31:0] T269;
  wire[31:0] T270;
  wire[31:0] T271;
  wire[31:0] T272;
  wire[31:0] T273;
  reg[31:0] linkIndex_1;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[31:0] T278;
  wire[31:0] T279;
  wire[31:0] T280;
  wire[31:0] T281;
  wire[31:0] T282;
  reg[31:0] linkIndex_0;
  wire T283;
  wire T284;
  wire T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire[31:0] T293;
  wire[31:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire[7:0] T299;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[31:0] T305;
  wire[31:0] T306;
  wire[31:0] T307;
  reg[31:0] pageId_0;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  reg[31:0] outPageId_1;
  wire[127:0] T319;
  wire[127:0] T320;
  wire[127:0] T321;
  wire[127:0] T322;
  wire[127:0] T323;
  reg[127:0] memRep_1_data;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[7:0] T330;
  wire T331;
  wire[127:0] T332;
  wire[127:0] T333;
  wire[127:0] T334;
  wire[127:0] T335;
  wire[127:0] T336;
  reg[127:0] memRep_0_data;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire[127:0] T342;
  wire[127:0] T343;
  wire[127:0] T344;
  wire[31:0] T345;
  wire[31:0] T346;
  reg[31:0] outPageId_0;
  wire[127:0] T347;
  wire[127:0] T348;
  wire[31:0] T349;
  wire[31:0] T350;
  reg[31:0] outputReg_0_pageId;
  wire T351;
  wire T352;
  wire[31:0] T353;
  wire[31:0] T354;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T355;
  wire[165:0] T356;
  wire[165:0] T357;
  wire[3:0] T358;
  wire[165:0] T359;
  wire[165:0] T360;
  wire[3:0] T361;
  wire[165:0] T362;
  wire[165:0] T363;
  wire[165:0] T364;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T365;
  wire[57:0] T366;
  wire[57:0] T367;
  wire[33:0] T368;
  wire[31:0] T369;
  wire[31:0] T370;
  wire[31:0] T371;
  reg[31:0] linkId_1;
  wire[127:0] T372;
  wire[127:0] T373;
  wire[127:0] T374;
  wire[31:0] T375;
  wire[31:0] T376;
  reg[31:0] linkId_0;
  wire[127:0] T377;
  wire[127:0] T378;
  wire T379;
  wire T380;
  wire[7:0] T381;
  wire T382;
  wire[127:0] T383;
  wire T384;
  wire T385;
  wire[31:0] T386;
  wire[165:0] T387;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T388;
  wire[34:0] T389;
  wire[34:0] T390;
  wire[31:0] T391;
  wire[31:0] T392;
  wire[31:0] T393;
  wire[31:0] T394;
  wire[31:0] T395;
  wire[34:0] T396;
  wire T397;
  wire T398;
  wire[7:0] T399;
  wire T400;
  wire[127:0] T401;
  wire T402;
  wire T403;
  wire[31:0] T404;
  wire[165:0] T405;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T406;
  wire[55:0] T407;
  wire[55:0] T408;
  wire[34:0] T409;
  wire T410;
  wire T411;
  wire[7:0] T412;
  wire T413;
  wire[127:0] T414;
  wire[127:0] T415;
  reg[127:0] memPortReplyStorage_0_data;
  wire T416;
  wire T417;
  wire[127:0] T418;
  wire[127:0] T419;
  wire T420;
  wire T421;
  wire[9:0] T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire[7:0] T442;
  wire[7:0] T443;
  wire[7:0] T444;
  wire[7:0] T445;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T448;
  wire[7:0] T449;
  wire[7:0] T450;
  wire[7:0] T451;
  wire[7:0] T452;
  wire[7:0] T453;
  wire[7:0] T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  reg[7:0] EmitReturnState_1;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  reg[7:0] EmitReturnState_0;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire[7:0] T514;
  wire[7:0] T515;
  wire[7:0] T516;
  wire[7:0] T517;
  wire[7:0] T518;
  wire[7:0] T519;
  wire[7:0] T520;
  wire[7:0] T521;
  wire[7:0] T522;
  wire[7:0] T523;
  wire[7:0] T524;
  wire[7:0] T525;
  wire[7:0] T526;
  wire[7:0] T527;
  wire[7:0] T528;
  wire[7:0] T529;
  wire[7:0] T530;
  wire[7:0] T531;
  wire[7:0] T532;
  wire[7:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire[1:0] T539;
  wire AllOffloadsReady;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  reg[0:0] rankCalcPortHadReadyRequest;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  reg[0:0] rankCalc_ready_received;
  wire T549;
  wire T550;
  wire rankCalcPort_req_ready;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  reg[0:0] memPortHadReadyRequest;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  reg[0:0] mem_ready_received;
  wire T560;
  wire T561;
  wire memPort_req_ready;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire T572;
  wire T573;
  wire[7:0] T574;
  wire[7:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[7:0] T580;
  wire T581;
  wire T582;
  wire T583;
  wire[7:0] T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T592;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T593;
  wire memPort_req_bits_cached;
  wire T594;
  wire memPort_req_bits_rw;
  wire T595;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T596;
  wire[9:0] T597;
  wire[9:0] T598;
  wire[9:0] T599;
  reg[9:0] inputTag_1;
  wire[9:0] T600;
  wire[9:0] T601;
  wire[9:0] T602;
  reg[9:0] inputTag_0;
  wire[9:0] T603;

  assign mainOff_mem_req_valid = memPort_req_valid;
  assign memPort_req_valid = T0;
  assign T0 = T586 && T1;
  assign T1 = T577 || T2;
  assign T2 = T576 && T3;
  assign T3 = T5 == T4;
  assign T4 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T5 = T574 | T6;
  assign T6 = State_1 & T7;
  assign T7 = {4'h8/* 8*/{T8}};
  assign T8 = T9[1'h1/* 1*/];
  assign T9 = T10[1'h1/* 1*/:1'h0/* 0*/];
  assign T10 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T11 = subStateTh_1 == 1'h0/* 0*/;
  assign T12 = T565 ? 1'h1/* 1*/ : T13;
  assign T13 = T14 ? 1'h0/* 0*/ : subStateTh_1;
  assign T14 = T564 == vThreadEncoder_io_chosen;
  assign T15 = T82 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T16;
  assign T16 = T60 && T17;
  assign T17 = T56 || T18;
  assign T18 = ! rankCalcPortHadValidRequest_1;
  assign T19 = T53 && T20;
  assign T20 = rankCalcPortHadValidRequest_1 || T21;
  assign T21 = T51 && rankCalcPort_req_valid;
  assign rankCalcPort_req_valid = T22;
  assign T22 = T27 && T23;
  assign T23 = T26 && T24;
  assign T24 = T5 == T25;
  assign T25 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T26 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T27 = T50 && T28;
  assign T28 = ! T29;
  assign T29 = T40 | T30;
  assign T30 = rankCalc_valid_received_1 & T8;
  assign T31 = T37 && T32;
  assign T32 = rankCalc_valid_received_1 || T33;
  assign T33 = rankCalcPort_rep_valid && T34;
  assign T34 = rankCalcPort_rep_tag == T35;
  assign T35 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign rankCalcPort_rep_tag = mainOff_rankCalc_rep_tag;
  assign mainOff_rankCalc_rep_ready = rankCalcPort_rep_ready;
  assign rankCalcPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_rankCalc_req_valid = rankCalcPort_req_valid;
  assign mainOff_rankCalc_req_tag = rankCalcPort_req_tag;
  assign rankCalcPort_req_tag = T36;
  assign T36 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign rankCalcPort_rep_valid = mainOff_rankCalc_rep_valid;
  assign T37 = ! T38;
  assign T38 = T39 == 5'h1/* 1*/;
  assign T39 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T40 = rankCalc_valid_received_0 & T41;
  assign T41 = T9[1'h0/* 0*/];
  assign T42 = T47 && T43;
  assign T43 = rankCalc_valid_received_0 || T44;
  assign T44 = rankCalcPort_rep_valid && T45;
  assign T45 = rankCalcPort_rep_tag == T46;
  assign T46 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T47 = ! T48;
  assign T48 = T49 == 5'h0/* 0*/;
  assign T49 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T50 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T51 = 5'h1/* 1*/ == T52;
  assign T52 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T53 = ! T54;
  assign T54 = T55 == 5'h1/* 1*/;
  assign T55 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T56 = T57 || rankCalc_valid_received_1;
  assign T57 = rankCalcPort_rep_valid && T58;
  assign T58 = rankCalcPort_rep_tag == T59;
  assign T59 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T60 = T70 || T61;
  assign T61 = ! memPortHadValidRequest_1;
  assign T62 = T67 && T63;
  assign T63 = memPortHadValidRequest_1 || T64;
  assign T64 = T65 && memPort_req_valid;
  assign T65 = 5'h1/* 1*/ == T66;
  assign T66 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T67 = ! T68;
  assign T68 = T69 == 5'h1/* 1*/;
  assign T69 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T70 = T79 || mem_valid_received_1;
  assign T71 = T76 && T72;
  assign T72 = mem_valid_received_1 || T73;
  assign T73 = memPort_rep_valid && T74;
  assign T74 = memPort_rep_tag == T75;
  assign T75 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T76 = ! T77;
  assign T77 = T78 == 5'h1/* 1*/;
  assign T78 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T79 = memPort_rep_valid && T80;
  assign T80 = memPort_rep_tag == T81;
  assign T81 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T82 = subStateTh_1 == 1'h1/* 1*/;
  assign T83 = T121 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T84;
  assign T84 = T99 && T85;
  assign T85 = T95 || T86;
  assign T86 = ! rankCalcPortHadValidRequest_0;
  assign T87 = T92 && T88;
  assign T88 = rankCalcPortHadValidRequest_0 || T89;
  assign T89 = T90 && rankCalcPort_req_valid;
  assign T90 = 5'h0/* 0*/ == T91;
  assign T91 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T92 = ! T93;
  assign T93 = T94 == 5'h0/* 0*/;
  assign T94 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T95 = T96 || rankCalc_valid_received_0;
  assign T96 = rankCalcPort_rep_valid && T97;
  assign T97 = rankCalcPort_rep_tag == T98;
  assign T98 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T99 = T109 || T100;
  assign T100 = ! memPortHadValidRequest_0;
  assign T101 = T106 && T102;
  assign T102 = memPortHadValidRequest_0 || T103;
  assign T103 = T104 && memPort_req_valid;
  assign T104 = 5'h0/* 0*/ == T105;
  assign T105 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T106 = ! T107;
  assign T107 = T108 == 5'h0/* 0*/;
  assign T108 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T109 = T118 || mem_valid_received_0;
  assign T110 = T115 && T111;
  assign T111 = mem_valid_received_0 || T112;
  assign T112 = memPort_rep_valid && T113;
  assign T113 = memPort_rep_tag == T114;
  assign T114 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T115 = ! T116;
  assign T116 = T117 == 5'h0/* 0*/;
  assign T117 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T118 = memPort_rep_valid && T119;
  assign T119 = memPort_rep_tag == T120;
  assign T120 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T121 = subStateTh_0 == 1'h1/* 1*/;
  assign T122 = T126 ? 1'h1/* 1*/ : T123;
  assign T123 = T124 ? 1'h0/* 0*/ : subStateTh_0;
  assign T124 = T125 == vThreadEncoder_io_chosen;
  assign T125 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T126 = T535 && T127;
  assign T127 = State_0 != 8'hff/* 255*/;
  assign T128 = T498 || T129;
  assign T129 = T133 && T130;
  assign T130 = T131[1'h0/* 0*/];
  assign T131 = T132[1'h1/* 1*/:1'h0/* 0*/];
  assign T132 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T133 = T497 && T134;
  assign T134 = T136 == T135;
  assign T135 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T136 = T495 | T137;
  assign T137 = State_1 & T138;
  assign T138 = {4'h8/* 8*/{T139}};
  assign T139 = T131[1'h1/* 1*/];
  assign T140 = T142 || T141;
  assign T141 = T133 && T139;
  assign T142 = T148 || T143;
  assign T143 = T144 && T139;
  assign T144 = T147 && T145;
  assign T145 = T136 == T146;
  assign T146 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T147 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T148 = T154 || T149;
  assign T149 = T150 && T139;
  assign T150 = T153 && T151;
  assign T151 = T136 == T152;
  assign T152 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T153 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T154 = T160 || T155;
  assign T155 = T156 && T139;
  assign T156 = T159 && T157;
  assign T157 = T136 == T158;
  assign T158 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T159 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T160 = T423 || T161;
  assign T161 = T162 && T139;
  assign T162 = T255 && T163;
  assign T163 = ! T164;
  assign T164 = page_fanoutDegree == 32'h0/* 0*/;
  assign page_fanoutDegree = T165;
  assign T165 = memRep1_data[5'h1f/* 31*/:1'h0/* 0*/];
  assign memRep1_data = T166;
  assign T166 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T420 ? T419 : T167;
  assign T167 = {T168};
  assign T168 = T414 | T169;
  assign T169 = memPortReplyStorage_1_data & T170;
  assign T170 = {8'h80/* 128*/{T139}};
  assign T171 = memPort_rep_valid && T172;
  assign T172 = T173[1'h1/* 1*/];
  assign T173 = T174[1'h1/* 1*/:1'h0/* 0*/];
  assign T174 = 2'h1/* 1*/ << memPort_rep_tag;
  assign T175 = T171 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign io_in_ready = T176;
  assign T176 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T177 = T179 && T178;
  assign T178 = State_1 == 8'h0/* 0*/;
  assign T179 = subStateTh_1 == 1'h0/* 0*/;
  assign T180 = T182 && T181;
  assign T181 = State_0 == 8'h0/* 0*/;
  assign T182 = subStateTh_0 == 1'h0/* 0*/;
  assign T183 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_valid = T184;
  assign T184 = T186 && T185;
  assign T185 = T5 == 8'hff/* 255*/;
  assign T186 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_bits_done = T187;
  assign T187 = T210 | T188;
  assign T188 = outputReg_1_done & T8;
  assign T189 = T190 || T141;
  assign T190 = T191 && T139;
  assign T191 = T194 && T192;
  assign T192 = T136 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T195 = T141 ? T197 : T196;
  assign T196 = T190 ? 1'h0/* 0*/ : outputReg_1_done;
  assign T197 = T206 | T198;
  assign T198 = inputReg_1_done & T139;
  assign T199 = T203 && T200;
  assign T200 = T201[1'h1/* 1*/];
  assign T201 = T202[1'h1/* 1*/:1'h0/* 0*/];
  assign T202 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T203 = T204 && io_in_valid;
  assign T204 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T205 = T199 ? io_in_bits_done : inputReg_1_done;
  assign T206 = inputReg_0_done & T130;
  assign T207 = T203 && T208;
  assign T208 = T201[1'h0/* 0*/];
  assign T209 = T207 ? io_in_bits_done : inputReg_0_done;
  assign T210 = outputReg_0_done & T41;
  assign T211 = T212 || T129;
  assign T212 = T191 && T130;
  assign T213 = T129 ? T197 : T214;
  assign T214 = T212 ? 1'h0/* 0*/ : outputReg_0_done;
  assign io_out_bits_pageId = T215;
  assign T215 = T349 | T216;
  assign T216 = outputReg_1_pageId & T217;
  assign T217 = {6'h20/* 32*/{T8}};
  assign T218 = T190 || T143;
  assign T219 = T143 ? T316 : T220;
  assign T220 = T190 ? T221 : outputReg_1_pageId;
  assign T221 = T306 | T222;
  assign T222 = pageId_1 & T223;
  assign T223 = {6'h20/* 32*/{T139}};
  assign T224 = T288 || T225;
  assign T225 = T226 && T139;
  assign T226 = T245 && T227;
  assign T227 = ! T228;
  assign T228 = T221 == T229;
  assign T229 = T230 - 32'h1/* 1*/;
  assign T230 = T238 + T231;
  assign T231 = T235 | T232;
  assign T232 = inputReg_1_length & T233;
  assign T233 = {6'h20/* 32*/{T139}};
  assign T234 = T199 ? io_in_bits_length : inputReg_1_length;
  assign T235 = inputReg_0_length & T236;
  assign T236 = {6'h20/* 32*/{T130}};
  assign T237 = T207 ? io_in_bits_length : inputReg_0_length;
  assign T238 = T242 | T239;
  assign T239 = inputReg_1_startPageId & T240;
  assign T240 = {6'h20/* 32*/{T139}};
  assign T241 = T199 ? io_in_bits_startPageId : inputReg_1_startPageId;
  assign T242 = inputReg_0_startPageId & T243;
  assign T243 = {6'h20/* 32*/{T130}};
  assign T244 = T207 ? io_in_bits_startPageId : inputReg_0_startPageId;
  assign T245 = T144 && T246;
  assign T246 = T271 == T247;
  assign T247 = T264 | T248;
  assign T248 = fanoutDegree_1 & T249;
  assign T249 = {6'h20/* 32*/{T139}};
  assign T250 = T259 || T251;
  assign T251 = T252 && T139;
  assign T252 = T255 && T253;
  assign T253 = ! T254;
  assign T254 = page_fanoutDegree <= 32'h20/* 32*/;
  assign T255 = T258 && T256;
  assign T256 = T136 == T257;
  assign T257 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T258 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T259 = T260 && T139;
  assign T260 = T255 && T254;
  assign T261 = T251 ? T263 : T262;
  assign T262 = T259 ? page_fanoutDegree : fanoutDegree_1;
  assign T263 = page_fanoutDegree & 32'h1f/* 31*/;
  assign T264 = fanoutDegree_0 & T265;
  assign T265 = {6'h20/* 32*/{T130}};
  assign T266 = T268 || T267;
  assign T267 = T252 && T130;
  assign T268 = T260 && T130;
  assign T269 = T267 ? T263 : T270;
  assign T270 = T268 ? page_fanoutDegree : fanoutDegree_0;
  assign T271 = T281 | T272;
  assign T272 = linkIndex_1 & T273;
  assign T273 = {6'h20/* 32*/{T139}};
  assign T274 = T155 || T275;
  assign T275 = T276 && T139;
  assign T276 = T144 && T277;
  assign T277 = ! T246;
  assign T278 = T275 ? T280 : T279;
  assign T279 = T155 ? 32'h0/* 0*/ : linkIndex_1;
  assign T280 = T271 + 32'h1/* 1*/;
  assign T281 = linkIndex_0 & T282;
  assign T282 = {6'h20/* 32*/{T130}};
  assign T283 = T285 || T284;
  assign T284 = T276 && T130;
  assign T285 = T156 && T130;
  assign T286 = T284 ? T280 : T287;
  assign T287 = T285 ? 32'h0/* 0*/ : linkIndex_0;
  assign T288 = T296 || T289;
  assign T289 = T290 && T139;
  assign T290 = T295 && T291;
  assign T291 = ! T292;
  assign T292 = T221 == T293;
  assign T293 = T294 - 32'h1/* 1*/;
  assign T294 = T238 + T231;
  assign T295 = T255 && T164;
  assign T296 = T297 && T139;
  assign T297 = T300 && T298;
  assign T298 = T136 == T299;
  assign T299 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T300 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T301 = T225 ? T305 : T302;
  assign T302 = T289 ? T304 : T303;
  assign T303 = T296 ? T238 : pageId_1;
  assign T304 = T221 + 32'h1/* 1*/;
  assign T305 = T221 + 32'h1/* 1*/;
  assign T306 = pageId_0 & T307;
  assign T307 = {6'h20/* 32*/{T130}};
  assign T308 = T310 || T309;
  assign T309 = T226 && T130;
  assign T310 = T312 || T311;
  assign T311 = T290 && T130;
  assign T312 = T297 && T130;
  assign T313 = T309 ? T305 : T314;
  assign T314 = T311 ? T304 : T315;
  assign T315 = T312 ? T238 : pageId_0;
  assign T316 = T345 | T317;
  assign T317 = outPageId_1 & T318;
  assign T318 = {6'h20/* 32*/{T139}};
  assign T319 = T149 ? T321 : T320;
  assign T320 = {96'h0/* 0*/, outPageId_1};
  assign T321 = T335 | T322;
  assign T322 = memRep_1_data & T323;
  assign T323 = {8'h80/* 128*/{T139}};
  assign T324 = T325 || T149;
  assign T325 = T327 || T326;
  assign T326 = T255 && T139;
  assign T327 = T328 && T139;
  assign T328 = T331 && T329;
  assign T329 = T136 == T330;
  assign T330 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T331 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T332 = T149 ? T166 : T333;
  assign T333 = T326 ? memRep1_data : T334;
  assign T334 = T327 ? T166 : memRep_1_data;
  assign T335 = memRep_0_data & T336;
  assign T336 = {8'h80/* 128*/{T130}};
  assign T337 = T339 || T338;
  assign T338 = T150 && T130;
  assign T339 = T341 || T340;
  assign T340 = T255 && T130;
  assign T341 = T328 && T130;
  assign T342 = T338 ? T166 : T343;
  assign T343 = T340 ? memRep1_data : T344;
  assign T344 = T341 ? T166 : memRep_0_data;
  assign T345 = outPageId_0 & T346;
  assign T346 = {6'h20/* 32*/{T130}};
  assign T347 = T338 ? T321 : T348;
  assign T348 = {96'h0/* 0*/, outPageId_0};
  assign T349 = outputReg_0_pageId & T350;
  assign T350 = {6'h20/* 32*/{T41}};
  assign T351 = T212 || T352;
  assign T352 = T144 && T130;
  assign T353 = T352 ? T316 : T354;
  assign T354 = T212 ? T221 : outputReg_0_pageId;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T355;
  assign T355 = T356[8'ha5/* 165*/:8'h86/* 134*/];
  assign T356 = T410 ? T405 : T357;
  assign T357 = {T404, T403, T402, T401, T358};
  assign T358 = T359[2'h3/* 3*/:1'h0/* 0*/];
  assign T359 = T397 ? T387 : T360;
  assign T360 = {T386, T385, T384, T383, T361};
  assign T361 = T362[2'h3/* 3*/:1'h0/* 0*/];
  assign T362 = T379 ? T364 : T363;
  assign T363 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T364 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h4/* 4*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T365;
  assign T365 = T366[5'h1f/* 31*/:1'h0/* 0*/];
  assign T366 = 58'h4000000/* 67108864*/ + T367;
  assign T367 = {24'h0/* 0*/, T368};
  assign T368 = T369 << 32'h2/* 2*/;
  assign T369 = T375 | T370;
  assign T370 = linkId_1 & T371;
  assign T371 = {6'h20/* 32*/{T8}};
  assign T372 = T326 ? T374 : T373;
  assign T373 = {96'h0/* 0*/, linkId_1};
  assign T374 = memRep1_data >> 32'h20/* 32*/;
  assign T375 = linkId_0 & T376;
  assign T376 = {6'h20/* 32*/{T41}};
  assign T377 = T340 ? T374 : T378;
  assign T378 = {96'h0/* 0*/, linkId_0};
  assign T379 = T382 && T380;
  assign T380 = T5 == T381;
  assign T381 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T382 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T383 = T362[8'h83/* 131*/:3'h4/* 4*/];
  assign T384 = T362[8'h84/* 132*/];
  assign T385 = T362[8'h85/* 133*/];
  assign T386 = T362[8'ha5/* 165*/:8'h86/* 134*/];
  assign T387 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h8/* 8*/;
  assign memReq2_cached = 1'h0/* 0*/;
  assign memReq2_rw = 1'h0/* 0*/;
  assign memReq2_addr = T388;
  assign T388 = T389[5'h1f/* 31*/:1'h0/* 0*/];
  assign T389 = T396 + T390;
  assign T390 = T391 << 32'h3/* 3*/;
  assign T391 = T394 | T392;
  assign T392 = pageId_1 & T393;
  assign T393 = {6'h20/* 32*/{T8}};
  assign T394 = pageId_0 & T395;
  assign T395 = {6'h20/* 32*/{T41}};
  assign T396 = {3'h0/* 0*/, 32'h0/* 0*/};
  assign T397 = T400 && T398;
  assign T398 = T5 == T399;
  assign T399 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T400 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T401 = T359[8'h83/* 131*/:3'h4/* 4*/];
  assign T402 = T359[8'h84/* 132*/];
  assign T403 = T359[8'h85/* 133*/];
  assign T404 = T359[8'ha5/* 165*/:8'h86/* 134*/];
  assign T405 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h8/* 8*/;
  assign memReq1_cached = 1'h0/* 0*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T406;
  assign T406 = T407[5'h1f/* 31*/:1'h0/* 0*/];
  assign T407 = 56'h1000000/* 16777216*/ + T408;
  assign T408 = {21'h0/* 0*/, T409};
  assign T409 = T391 << 32'h3/* 3*/;
  assign T410 = T413 && T411;
  assign T411 = T5 == T412;
  assign T412 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T413 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T414 = memPortReplyStorage_0_data & T415;
  assign T415 = {8'h80/* 128*/{T130}};
  assign T416 = memPort_rep_valid && T417;
  assign T417 = T173[1'h0/* 0*/];
  assign T418 = T416 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T419 = {memPort_rep_bits_data};
  assign T420 = memPort_rep_valid && T421;
  assign T421 = T422 == memPort_rep_tag;
  assign T422 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T423 = T424 || T289;
  assign T424 = T427 || T425;
  assign T425 = T426 && T139;
  assign T426 = T295 && T292;
  assign T427 = T428 || T327;
  assign T428 = T429 || T190;
  assign T429 = T433 || T430;
  assign T430 = T431 && T139;
  assign T431 = T297 && T432;
  assign T432 = ! T197;
  assign T433 = T436 || T434;
  assign T434 = T435 && T139;
  assign T435 = T297 && T197;
  assign T436 = T199 || T437;
  assign T437 = T438 && T8;
  assign T438 = T439 && io_out_ready;
  assign T439 = T441 && T440;
  assign T440 = T5 == 8'hff/* 255*/;
  assign T441 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T442 = T494 ? 8'hff/* 255*/ : T443;
  assign T443 = T149 ? T493 : T444;
  assign T444 = T155 ? T492 : T445;
  assign T445 = T161 ? T491 : T446;
  assign T446 = T289 ? T490 : T447;
  assign T447 = T425 ? 8'h0/* 0*/ : T448;
  assign T448 = T327 ? T489 : T449;
  assign T449 = T190 ? 8'hff/* 255*/ : T450;
  assign T450 = T430 ? T488 : T451;
  assign T451 = T434 ? T487 : T452;
  assign T452 = T437 ? T455 : T453;
  assign T453 = T199 ? T454 : State_1;
  assign T454 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T455 = T472 | T456;
  assign T456 = EmitReturnState_1 & T457;
  assign T457 = {4'h8/* 8*/{T8}};
  assign T458 = T459 || T141;
  assign T459 = T460 || T275;
  assign T460 = T461 || T225;
  assign T461 = T190 || T462;
  assign T462 = T463 && T139;
  assign T463 = T245 && T228;
  assign T464 = T141 ? 8'h0/* 0*/ : T465;
  assign T465 = T275 ? T471 : T466;
  assign T466 = T225 ? T470 : T467;
  assign T467 = T462 ? 8'h0/* 0*/ : T468;
  assign T468 = T190 ? T469 : EmitReturnState_1;
  assign T469 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T470 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T471 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T472 = EmitReturnState_0 & T473;
  assign T473 = {4'h8/* 8*/{T41}};
  assign T474 = T475 || T129;
  assign T475 = T476 || T284;
  assign T476 = T477 || T309;
  assign T477 = T212 || T478;
  assign T478 = T463 && T130;
  assign T479 = T129 ? 8'h0/* 0*/ : T480;
  assign T480 = T284 ? T486 : T481;
  assign T481 = T309 ? T485 : T482;
  assign T482 = T478 ? 8'h0/* 0*/ : T483;
  assign T483 = T212 ? T484 : EmitReturnState_0;
  assign T484 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T485 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T486 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T487 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T488 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T489 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T492 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T493 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T494 = T143 || T141;
  assign T495 = State_0 & T496;
  assign T496 = {4'h8/* 8*/{T130}};
  assign T497 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T498 = T499 || T352;
  assign T499 = T500 || T338;
  assign T500 = T501 || T285;
  assign T501 = T503 || T502;
  assign T502 = T162 && T130;
  assign T503 = T504 || T311;
  assign T504 = T506 || T505;
  assign T505 = T426 && T130;
  assign T506 = T507 || T341;
  assign T507 = T508 || T212;
  assign T508 = T510 || T509;
  assign T509 = T431 && T130;
  assign T510 = T512 || T511;
  assign T511 = T435 && T130;
  assign T512 = T207 || T513;
  assign T513 = T438 && T41;
  assign T514 = T534 ? 8'hff/* 255*/ : T515;
  assign T515 = T338 ? T533 : T516;
  assign T516 = T285 ? T532 : T517;
  assign T517 = T502 ? T531 : T518;
  assign T518 = T311 ? T530 : T519;
  assign T519 = T505 ? 8'h0/* 0*/ : T520;
  assign T520 = T341 ? T529 : T521;
  assign T521 = T212 ? 8'hff/* 255*/ : T522;
  assign T522 = T509 ? T528 : T523;
  assign T523 = T511 ? T527 : T524;
  assign T524 = T513 ? T455 : T525;
  assign T525 = T207 ? T526 : State_0;
  assign T526 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T527 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T528 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T529 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T530 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T531 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T532 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T533 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T534 = T352 || T129;
  assign T535 = T537 && T536;
  assign T536 = State_0 != 8'h0/* 0*/;
  assign T537 = AllOffloadsReady && T538;
  assign T538 = T539 == rThreadEncoder_io_chosen;
  assign T539 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign AllOffloadsReady = T540;
  assign T540 = T552 && T541;
  assign T541 = T548 || T542;
  assign T542 = T544 && T543;
  assign T543 = ! rankCalcPort_req_valid;
  assign T544 = ! rankCalcPortHadReadyRequest;
  assign T545 = T547 && T546;
  assign T546 = rankCalcPortHadReadyRequest || rankCalcPort_req_valid;
  assign T547 = ! AllOffloadsReady;
  assign T548 = rankCalcPort_req_ready || rankCalc_ready_received;
  assign T549 = T551 && T550;
  assign T550 = rankCalc_ready_received || rankCalcPort_req_ready;
  assign rankCalcPort_req_ready = mainOff_rankCalc_req_ready;
  assign T551 = ! AllOffloadsReady;
  assign T552 = T559 || T553;
  assign T553 = T555 && T554;
  assign T554 = ! memPort_req_valid;
  assign T555 = ! memPortHadReadyRequest;
  assign T556 = T558 && T557;
  assign T557 = memPortHadReadyRequest || memPort_req_valid;
  assign T558 = ! AllOffloadsReady;
  assign T559 = memPort_req_ready || mem_ready_received;
  assign T560 = T562 && T561;
  assign T561 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign T562 = ! AllOffloadsReady;
  assign T563 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T564 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T565 = T567 && T566;
  assign T566 = State_1 != 8'hff/* 255*/;
  assign T567 = T569 && T568;
  assign T568 = State_1 != 8'h0/* 0*/;
  assign T569 = AllOffloadsReady && T570;
  assign T570 = T571 == rThreadEncoder_io_chosen;
  assign T571 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T572 = subStateTh_0 == 1'h0/* 0*/;
  assign T573 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T574 = State_0 & T575;
  assign T575 = {4'h8/* 8*/{T41}};
  assign T576 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T577 = T582 || T578;
  assign T578 = T581 && T579;
  assign T579 = T5 == T580;
  assign T580 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T581 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T582 = T585 && T583;
  assign T583 = T5 == T584;
  assign T584 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T585 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T586 = T591 && T587;
  assign T587 = ! T588;
  assign T588 = T590 | T589;
  assign T589 = mem_valid_received_1 & T8;
  assign T590 = mem_valid_received_0 & T41;
  assign T591 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T592;
  assign T592 = T356[2'h3/* 3*/:1'h0/* 0*/];
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T593;
  assign T593 = T356[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T594;
  assign T594 = T356[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T595;
  assign T595 = T356[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T596;
  assign T596 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign io_out_tag = T597;
  assign T597 = T601 | T598;
  assign T598 = inputTag_1 & T599;
  assign T599 = {4'ha/* 10*/{T8}};
  assign T600 = T199 ? io_in_tag : inputTag_1;
  assign T601 = inputTag_0 & T602;
  assign T602 = {4'ha/* 10*/{T41}};
  assign T603 = T207 ? io_in_tag : inputTag_0;
  RREncode rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T572 ),
       .io_valid_1( T11 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T573 ));
  RREncode_1 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T83 ),
       .io_valid_1( T15 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T563 ));
  RREncode_2 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T180 ),
       .io_valid_1( T177 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T183 ));

  always @(posedge clk) begin
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T12;
    rankCalcPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T19;
    rankCalc_valid_received_1 <= reset ? 1'h0/* 0*/ : T31;
    rankCalc_valid_received_0 <= reset ? 1'h0/* 0*/ : T42;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T62;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T71;
    rankCalcPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T87;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T101;
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T110;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T122;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T128) begin
      State_0 <= T514;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T140) begin
      State_1 <= T442;
    end
    if(T171) begin
      memPortReplyStorage_1_data <= T175;
    end
    if(T189) begin
      outputReg_1_done <= T195;
    end
    if(T199) begin
      inputReg_1_done <= T205;
    end
    if(T207) begin
      inputReg_0_done <= T209;
    end
    if(T211) begin
      outputReg_0_done <= T213;
    end
    if(T218) begin
      outputReg_1_pageId <= T219;
    end
    if(T224) begin
      pageId_1 <= T301;
    end
    if(T199) begin
      inputReg_1_length <= T234;
    end
    if(T207) begin
      inputReg_0_length <= T237;
    end
    if(T199) begin
      inputReg_1_startPageId <= T241;
    end
    if(T207) begin
      inputReg_0_startPageId <= T244;
    end
    if(T250) begin
      fanoutDegree_1 <= T261;
    end
    if(T266) begin
      fanoutDegree_0 <= T269;
    end
    if(T274) begin
      linkIndex_1 <= T278;
    end
    if(T283) begin
      linkIndex_0 <= T286;
    end
    if(T308) begin
      pageId_0 <= T313;
    end
    if(T149) begin
      outPageId_1 <= T319;
    end
    if(T324) begin
      memRep_1_data <= T332;
    end
    if(T337) begin
      memRep_0_data <= T342;
    end
    if(T338) begin
      outPageId_0 <= T347;
    end
    if(T351) begin
      outputReg_0_pageId <= T353;
    end
    if(T326) begin
      linkId_1 <= T372;
    end
    if(T340) begin
      linkId_0 <= T377;
    end
    if(T416) begin
      memPortReplyStorage_0_data <= T418;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T458) begin
      EmitReturnState_1 <= T464;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T474) begin
      EmitReturnState_0 <= T479;
    end
    rankCalcPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T545;
    rankCalc_ready_received <= reset ? 1'h0/* 0*/ : T549;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T556;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T560;
    if(T199) begin
      inputTag_1 <= T600;
    end
    if(T207) begin
      inputTag_0 <= T603;
    end
  end
endmodule

module RREncode_3(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_4(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_5(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_6(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module rankCalculator(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  outputReg_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mul_req_ready,
    output mainOff_mul_req_valid,
    output[63:0] mainOff_mul_req_bits_in1,
    output[63:0] mainOff_mul_req_bits_in2,
    output[9:0] mainOff_mul_req_tag,
    output mainOff_mul_rep_ready,
    input  mainOff_mul_rep_valid,
    input [63:0] mainOff_mul_rep_bits_out,
    input [9:0] mainOff_mul_rep_tag,
    input  mainOff_div_req_ready,
    output mainOff_div_req_valid,
    output[63:0] mainOff_div_req_bits_in1,
    output[63:0] mainOff_div_req_bits_in2,
    output[9:0] mainOff_div_req_tag,
    output mainOff_div_rep_ready,
    input  mainOff_div_rep_valid,
    input [63:0] mainOff_div_rep_bits_out,
    input [9:0] mainOff_div_rep_tag);

  reg[9:0] outputReg_tag;
  wire T0;
  wire T1;
  wire[2:0] GS_step2VThreadEncoder_io_chosen;
  wire T2;
  wire GS_step2AllOffloadsValid_3;
  wire T3;
  wire T4;
  reg[0:0] mulPortHadValidRequest_3;
  wire T5;
  wire T6;
  wire T7;
  wire mulPort_req_valid;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] GS_step2RThreadEncoder_io_chosen;
  wire T11;
  reg[0:0] GS_step2PRegPostOff_valid_3;
  wire T12;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire[10:0] T16;
  wire GS_step2PipeValidMove;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire GS_step2AllOffloadsValid_2;
  wire T23;
  wire T24;
  reg[0:0] mulPortHadValidRequest_2;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[9:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire[9:0] T33;
  wire T34;
  reg[0:0] mulValidReceived_2;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[9:0] mulPort_rep_tag;
  wire mulPort_rep_ready;
  wire[9:0] mulPort_req_tag;
  wire[9:0] T39;
  wire mulPort_rep_valid;
  wire T40;
  wire T41;
  wire T42;
  wire[9:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire GS_step2AllOffloadsValid_1;
  wire T49;
  wire T50;
  reg[0:0] mulPortHadValidRequest_1;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[9:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[9:0] T59;
  wire T60;
  reg[0:0] mulValidReceived_1;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[9:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire GS_step2AllOffloadsValid_0;
  wire T73;
  wire T74;
  reg[0:0] mulPortHadValidRequest_0;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire[9:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire[9:0] T83;
  wire T84;
  reg[0:0] mulValidReceived_0;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[3:0] T99;
  wire[10:0] T100;
  wire T101;
  wire GS_step2AllOffloadsReady;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  reg[0:0] mulPortHadReadyRequest;
  wire T106;
  wire T107;
  wire T108;
  wire GS_step2PipeReadyMove;
  wire T109;
  wire T110;
  wire GS_step2PRegPostOff_ready;
  wire T111;
  wire T112;
  wire T113;
  reg[0:0] mulReadyReceived;
  wire T114;
  wire T115;
  wire mulPort_req_ready;
  wire T116;
  wire T117;
  reg[0:0] GS_step2PRegPreOff_valid;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] GS_step1VThreadEncoder_io_chosen;
  wire T122;
  wire GS_step1AllOffloadsValid_3;
  wire T123;
  wire T124;
  reg[0:0] divPortHadValidRequest_3;
  wire T125;
  wire T126;
  wire T127;
  wire divPort_req_valid;
  wire T128;
  wire T129;
  wire T130;
  wire[2:0] GS_step1RThreadEncoder_io_chosen;
  wire T131;
  reg[0:0] GS_step1PRegPostOff_valid_3;
  wire T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire[10:0] T136;
  wire GS_step1PipeValidMove;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire GS_step1AllOffloadsValid_2;
  wire T143;
  wire T144;
  reg[0:0] divPortHadValidRequest_2;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire[9:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire[9:0] T153;
  wire T154;
  reg[0:0] divValidReceived_2;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[9:0] divPort_rep_tag;
  wire divPort_rep_ready;
  wire[9:0] divPort_req_tag;
  wire[9:0] T159;
  wire divPort_rep_valid;
  wire T160;
  wire T161;
  wire T162;
  wire[9:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire GS_step1AllOffloadsValid_1;
  wire T169;
  wire T170;
  reg[0:0] divPortHadValidRequest_1;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[9:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire[9:0] T179;
  wire T180;
  reg[0:0] divValidReceived_1;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[9:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire GS_step1AllOffloadsValid_0;
  wire T193;
  wire T194;
  reg[0:0] divPortHadValidRequest_0;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire[9:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire[9:0] T203;
  wire T204;
  reg[0:0] divValidReceived_0;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[9:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire GS_step2PRegPreOff_ready;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[3:0] T220;
  wire[10:0] T221;
  wire T222;
  wire GS_step1AllOffloadsReady;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  reg[0:0] divPortHadReadyRequest;
  wire T227;
  wire T228;
  wire T229;
  wire GS_step1PipeReadyMove;
  wire T230;
  wire T231;
  wire GS_step1PRegPostOff_ready;
  wire T232;
  wire T233;
  wire T234;
  reg[0:0] divReadyReceived;
  wire T235;
  wire T236;
  wire divPort_req_ready;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  reg[0:0] GS_step1PRegPostOff_valid_2;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  reg[0:0] GS_step1PRegPostOff_valid_1;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  reg[0:0] GS_step1PRegPostOff_valid_0;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  reg[0:0] divValidReceived_3;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire[9:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[9:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire[9:0] T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  reg[0:0] GS_step2PRegPostOff_valid_2;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  reg[0:0] GS_step2PRegPostOff_valid_1;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  reg[0:0] GS_step2PRegPostOff_valid_0;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] mulValidReceived_3;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire[9:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire[9:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire[9:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  reg[0:0] outputReg_valid;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[9:0] T370;
  wire[9:0] T371;
  wire[9:0] T372;
  wire[9:0] T373;
  wire[9:0] T374;
  reg[9:0] GS_step2PRegPostOff_tag_3;
  wire[9:0] T375;
  wire[9:0] T376;
  reg[9:0] GS_step2PRegPreOff_tag;
  wire[9:0] T377;
  wire[9:0] T378;
  wire[9:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  reg[9:0] GS_step1PRegPostOff_tag_3;
  wire[9:0] T382;
  wire[9:0] T383;
  wire[9:0] T384;
  wire[9:0] T385;
  wire[9:0] T386;
  reg[9:0] GS_step1PRegPostOff_tag_2;
  wire[9:0] T387;
  wire[9:0] T388;
  wire[9:0] T389;
  wire[9:0] T390;
  wire[9:0] T391;
  reg[9:0] GS_step1PRegPostOff_tag_1;
  wire[9:0] T392;
  wire[9:0] T393;
  wire[9:0] T394;
  wire[9:0] T395;
  reg[9:0] GS_step1PRegPostOff_tag_0;
  wire[9:0] T396;
  wire[9:0] T397;
  wire[9:0] T398;
  wire[9:0] T399;
  wire[9:0] T400;
  reg[9:0] GS_step2PRegPostOff_tag_2;
  wire[9:0] T401;
  wire[9:0] T402;
  wire[9:0] T403;
  wire[9:0] T404;
  wire[9:0] T405;
  reg[9:0] GS_step2PRegPostOff_tag_1;
  wire[9:0] T406;
  wire[9:0] T407;
  wire[9:0] T408;
  wire[9:0] T409;
  reg[9:0] GS_step2PRegPostOff_tag_0;
  wire[9:0] T410;
  wire[9:0] T411;
  wire T412;

  assign io_out_tag = outputReg_tag;
  assign T0 = T356 && T1;
  assign T1 = GS_step2VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T2 = GS_step2PRegPostOff_valid_3 && GS_step2AllOffloadsValid_3;
  assign GS_step2AllOffloadsValid_3 = T3;
  assign T3 = T350 || T4;
  assign T4 = ! mulPortHadValidRequest_3;
  assign T5 = T346 && T6;
  assign T6 = mulPortHadValidRequest_3 || T7;
  assign T7 = T344 && mulPort_req_valid;
  assign mulPort_req_valid = T8;
  assign T8 = T326 && T9;
  assign T9 = GS_step2PRegPreOff_valid && T10;
  assign T10 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T11 = ! GS_step2PRegPostOff_valid_3;
  assign T12 = T97 || T13;
  assign T13 = GS_step2PipeValidMove && T14;
  assign T14 = T15[2'h3/* 3*/];
  assign T15 = T16[2'h3/* 3*/:1'h0/* 0*/];
  assign T16 = 4'h1/* 1*/ << GS_step2VThreadEncoder_io_chosen;
  assign GS_step2PipeValidMove = T17;
  assign T17 = T95 && T18;
  assign T18 = T20 | T19;
  assign T19 = GS_step2AllOffloadsValid_3 & T14;
  assign T20 = T46 | T21;
  assign T21 = GS_step2AllOffloadsValid_2 & T22;
  assign T22 = T15[2'h2/* 2*/];
  assign GS_step2AllOffloadsValid_2 = T23;
  assign T23 = T34 || T24;
  assign T24 = ! mulPortHadValidRequest_2;
  assign T25 = T30 && T26;
  assign T26 = mulPortHadValidRequest_2 || T27;
  assign T27 = T28 && mulPort_req_valid;
  assign T28 = 10'h2/* 2*/ == T29;
  assign T29 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T30 = ! T31;
  assign T31 = GS_step2PipeValidMove && T32;
  assign T32 = T33 == 10'h2/* 2*/;
  assign T33 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T34 = T44 || mulValidReceived_2;
  assign T35 = T40 && T36;
  assign T36 = mulValidReceived_2 || T37;
  assign T37 = mulPort_rep_valid && T38;
  assign T38 = mulPort_rep_tag == 10'h2/* 2*/;
  assign mulPort_rep_tag = mainOff_mul_rep_tag;
  assign mainOff_mul_rep_ready = mulPort_rep_ready;
  assign mulPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul_req_tag = mulPort_req_tag;
  assign mulPort_req_tag = T39;
  assign T39 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign mulPort_rep_valid = mainOff_mul_rep_valid;
  assign mainOff_mul_req_valid = mulPort_req_valid;
  assign T40 = ! T41;
  assign T41 = GS_step2PipeValidMove && T42;
  assign T42 = T43 == 10'h2/* 2*/;
  assign T43 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T44 = mulPort_rep_valid && T45;
  assign T45 = mulPort_rep_tag == 10'h2/* 2*/;
  assign T46 = T71 | T47;
  assign T47 = GS_step2AllOffloadsValid_1 & T48;
  assign T48 = T15[1'h1/* 1*/];
  assign GS_step2AllOffloadsValid_1 = T49;
  assign T49 = T60 || T50;
  assign T50 = ! mulPortHadValidRequest_1;
  assign T51 = T56 && T52;
  assign T52 = mulPortHadValidRequest_1 || T53;
  assign T53 = T54 && mulPort_req_valid;
  assign T54 = 10'h1/* 1*/ == T55;
  assign T55 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T56 = ! T57;
  assign T57 = GS_step2PipeValidMove && T58;
  assign T58 = T59 == 10'h1/* 1*/;
  assign T59 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T60 = T69 || mulValidReceived_1;
  assign T61 = T65 && T62;
  assign T62 = mulValidReceived_1 || T63;
  assign T63 = mulPort_rep_valid && T64;
  assign T64 = mulPort_rep_tag == 10'h1/* 1*/;
  assign T65 = ! T66;
  assign T66 = GS_step2PipeValidMove && T67;
  assign T67 = T68 == 10'h1/* 1*/;
  assign T68 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T69 = mulPort_rep_valid && T70;
  assign T70 = mulPort_rep_tag == 10'h1/* 1*/;
  assign T71 = GS_step2AllOffloadsValid_0 & T72;
  assign T72 = T15[1'h0/* 0*/];
  assign GS_step2AllOffloadsValid_0 = T73;
  assign T73 = T84 || T74;
  assign T74 = ! mulPortHadValidRequest_0;
  assign T75 = T80 && T76;
  assign T76 = mulPortHadValidRequest_0 || T77;
  assign T77 = T78 && mulPort_req_valid;
  assign T78 = 10'h0/* 0*/ == T79;
  assign T79 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T80 = ! T81;
  assign T81 = GS_step2PipeValidMove && T82;
  assign T82 = T83 == 10'h0/* 0*/;
  assign T83 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T84 = T93 || mulValidReceived_0;
  assign T85 = T89 && T86;
  assign T86 = mulValidReceived_0 || T87;
  assign T87 = mulPort_rep_valid && T88;
  assign T88 = mulPort_rep_tag == 10'h0/* 0*/;
  assign T89 = ! T90;
  assign T90 = GS_step2PipeValidMove && T91;
  assign T91 = T92 == 10'h0/* 0*/;
  assign T92 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T93 = mulPort_rep_valid && T94;
  assign T94 = mulPort_rep_tag == 10'h0/* 0*/;
  assign T95 = T96 && outputReg_ready;
  assign T96 = GS_step2VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T97 = T101 && T98;
  assign T98 = T99[2'h3/* 3*/];
  assign T99 = T100[2'h3/* 3*/:1'h0/* 0*/];
  assign T100 = 4'h1/* 1*/ << GS_step2RThreadEncoder_io_chosen;
  assign T101 = T117 && GS_step2AllOffloadsReady;
  assign GS_step2AllOffloadsReady = T102;
  assign T102 = T113 || T103;
  assign T103 = T105 && T104;
  assign T104 = ! mulPort_req_valid;
  assign T105 = ! mulPortHadReadyRequest;
  assign T106 = T108 && T107;
  assign T107 = mulPortHadReadyRequest || mulPort_req_valid;
  assign T108 = ! GS_step2PipeReadyMove;
  assign GS_step2PipeReadyMove = T109;
  assign T109 = T110 && GS_step2AllOffloadsReady;
  assign T110 = T112 && GS_step2PRegPostOff_ready;
  assign GS_step2PRegPostOff_ready = T111;
  assign T111 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T112 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T113 = mulPort_req_ready || mulReadyReceived;
  assign T114 = T116 && T115;
  assign T115 = mulReadyReceived || mulPort_req_ready;
  assign mulPort_req_ready = mainOff_mul_req_ready;
  assign T116 = ! GS_step2PipeReadyMove;
  assign T117 = GS_step2PRegPreOff_valid && GS_step2PRegPostOff_ready;
  assign T118 = T293 || T119;
  assign T119 = T291 && T120;
  assign T120 = ! T121;
  assign T121 = GS_step1VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T122 = GS_step1PRegPostOff_valid_3 && GS_step1AllOffloadsValid_3;
  assign GS_step1AllOffloadsValid_3 = T123;
  assign T123 = T285 || T124;
  assign T124 = ! divPortHadValidRequest_3;
  assign T125 = T281 && T126;
  assign T126 = divPortHadValidRequest_3 || T127;
  assign T127 = T279 && divPort_req_valid;
  assign divPort_req_valid = T128;
  assign T128 = T261 && T129;
  assign T129 = io_in_valid && T130;
  assign T130 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T131 = ! GS_step1PRegPostOff_valid_3;
  assign T132 = T218 || T133;
  assign T133 = GS_step1PipeValidMove && T134;
  assign T134 = T135[2'h3/* 3*/];
  assign T135 = T136[2'h3/* 3*/:1'h0/* 0*/];
  assign T136 = 4'h1/* 1*/ << GS_step1VThreadEncoder_io_chosen;
  assign GS_step1PipeValidMove = T137;
  assign T137 = T215 && T138;
  assign T138 = T140 | T139;
  assign T139 = GS_step1AllOffloadsValid_3 & T134;
  assign T140 = T166 | T141;
  assign T141 = GS_step1AllOffloadsValid_2 & T142;
  assign T142 = T135[2'h2/* 2*/];
  assign GS_step1AllOffloadsValid_2 = T143;
  assign T143 = T154 || T144;
  assign T144 = ! divPortHadValidRequest_2;
  assign T145 = T150 && T146;
  assign T146 = divPortHadValidRequest_2 || T147;
  assign T147 = T148 && divPort_req_valid;
  assign T148 = 10'h2/* 2*/ == T149;
  assign T149 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T150 = ! T151;
  assign T151 = GS_step1PipeValidMove && T152;
  assign T152 = T153 == 10'h2/* 2*/;
  assign T153 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T154 = T164 || divValidReceived_2;
  assign T155 = T160 && T156;
  assign T156 = divValidReceived_2 || T157;
  assign T157 = divPort_rep_valid && T158;
  assign T158 = divPort_rep_tag == 10'h2/* 2*/;
  assign divPort_rep_tag = mainOff_div_rep_tag;
  assign mainOff_div_rep_ready = divPort_rep_ready;
  assign divPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_div_req_tag = divPort_req_tag;
  assign divPort_req_tag = T159;
  assign T159 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign divPort_rep_valid = mainOff_div_rep_valid;
  assign mainOff_div_req_valid = divPort_req_valid;
  assign T160 = ! T161;
  assign T161 = GS_step1PipeValidMove && T162;
  assign T162 = T163 == 10'h2/* 2*/;
  assign T163 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T164 = divPort_rep_valid && T165;
  assign T165 = divPort_rep_tag == 10'h2/* 2*/;
  assign T166 = T191 | T167;
  assign T167 = GS_step1AllOffloadsValid_1 & T168;
  assign T168 = T135[1'h1/* 1*/];
  assign GS_step1AllOffloadsValid_1 = T169;
  assign T169 = T180 || T170;
  assign T170 = ! divPortHadValidRequest_1;
  assign T171 = T176 && T172;
  assign T172 = divPortHadValidRequest_1 || T173;
  assign T173 = T174 && divPort_req_valid;
  assign T174 = 10'h1/* 1*/ == T175;
  assign T175 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T176 = ! T177;
  assign T177 = GS_step1PipeValidMove && T178;
  assign T178 = T179 == 10'h1/* 1*/;
  assign T179 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T180 = T189 || divValidReceived_1;
  assign T181 = T185 && T182;
  assign T182 = divValidReceived_1 || T183;
  assign T183 = divPort_rep_valid && T184;
  assign T184 = divPort_rep_tag == 10'h1/* 1*/;
  assign T185 = ! T186;
  assign T186 = GS_step1PipeValidMove && T187;
  assign T187 = T188 == 10'h1/* 1*/;
  assign T188 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T189 = divPort_rep_valid && T190;
  assign T190 = divPort_rep_tag == 10'h1/* 1*/;
  assign T191 = GS_step1AllOffloadsValid_0 & T192;
  assign T192 = T135[1'h0/* 0*/];
  assign GS_step1AllOffloadsValid_0 = T193;
  assign T193 = T204 || T194;
  assign T194 = ! divPortHadValidRequest_0;
  assign T195 = T200 && T196;
  assign T196 = divPortHadValidRequest_0 || T197;
  assign T197 = T198 && divPort_req_valid;
  assign T198 = 10'h0/* 0*/ == T199;
  assign T199 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T200 = ! T201;
  assign T201 = GS_step1PipeValidMove && T202;
  assign T202 = T203 == 10'h0/* 0*/;
  assign T203 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T204 = T213 || divValidReceived_0;
  assign T205 = T209 && T206;
  assign T206 = divValidReceived_0 || T207;
  assign T207 = divPort_rep_valid && T208;
  assign T208 = divPort_rep_tag == 10'h0/* 0*/;
  assign T209 = ! T210;
  assign T210 = GS_step1PipeValidMove && T211;
  assign T211 = T212 == 10'h0/* 0*/;
  assign T212 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T213 = divPort_rep_valid && T214;
  assign T214 = divPort_rep_tag == 10'h0/* 0*/;
  assign T215 = T217 && GS_step2PRegPreOff_ready;
  assign GS_step2PRegPreOff_ready = T216;
  assign T216 = GS_step2PRegPostOff_ready && GS_step2AllOffloadsReady;
  assign T217 = GS_step1VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T218 = T222 && T219;
  assign T219 = T220[2'h3/* 3*/];
  assign T220 = T221[2'h3/* 3*/:1'h0/* 0*/];
  assign T221 = 4'h1/* 1*/ << GS_step1RThreadEncoder_io_chosen;
  assign T222 = GS_step1PRegPostOff_ready && GS_step1AllOffloadsReady;
  assign GS_step1AllOffloadsReady = T223;
  assign T223 = T234 || T224;
  assign T224 = T226 && T225;
  assign T225 = ! divPort_req_valid;
  assign T226 = ! divPortHadReadyRequest;
  assign T227 = T229 && T228;
  assign T228 = divPortHadReadyRequest || divPort_req_valid;
  assign T229 = ! GS_step1PipeReadyMove;
  assign GS_step1PipeReadyMove = T230;
  assign T230 = T231 && GS_step1AllOffloadsReady;
  assign T231 = T233 && GS_step1PRegPostOff_ready;
  assign GS_step1PRegPostOff_ready = T232;
  assign T232 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T233 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T234 = divPort_req_ready || divReadyReceived;
  assign T235 = T237 && T236;
  assign T236 = divReadyReceived || divPort_req_ready;
  assign divPort_req_ready = mainOff_div_req_ready;
  assign T237 = ! GS_step1PipeReadyMove;
  assign T238 = T133 ? 1'h0/* 0*/ : T239;
  assign T239 = T218 ? io_in_valid : GS_step1PRegPostOff_valid_3;
  assign T240 = ! GS_step1PRegPostOff_valid_2;
  assign T241 = T243 || T242;
  assign T242 = GS_step1PipeValidMove && T142;
  assign T243 = T222 && T244;
  assign T244 = T220[2'h2/* 2*/];
  assign T245 = T242 ? 1'h0/* 0*/ : T246;
  assign T246 = T243 ? io_in_valid : GS_step1PRegPostOff_valid_2;
  assign T247 = ! GS_step1PRegPostOff_valid_1;
  assign T248 = T250 || T249;
  assign T249 = GS_step1PipeValidMove && T168;
  assign T250 = T222 && T251;
  assign T251 = T220[1'h1/* 1*/];
  assign T252 = T249 ? 1'h0/* 0*/ : T253;
  assign T253 = T250 ? io_in_valid : GS_step1PRegPostOff_valid_1;
  assign T254 = ! GS_step1PRegPostOff_valid_0;
  assign T255 = T257 || T256;
  assign T256 = GS_step1PipeValidMove && T192;
  assign T257 = T222 && T258;
  assign T258 = T220[1'h0/* 0*/];
  assign T259 = T256 ? 1'h0/* 0*/ : T260;
  assign T260 = T257 ? io_in_valid : GS_step1PRegPostOff_valid_0;
  assign T261 = T278 && T262;
  assign T262 = ! T263;
  assign T263 = T273 | T264;
  assign T264 = divValidReceived_3 & T219;
  assign T265 = T269 && T266;
  assign T266 = divValidReceived_3 || T267;
  assign T267 = divPort_rep_valid && T268;
  assign T268 = divPort_rep_tag == 10'h3/* 3*/;
  assign T269 = ! T270;
  assign T270 = GS_step1PipeValidMove && T271;
  assign T271 = T272 == 10'h3/* 3*/;
  assign T272 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T273 = T275 | T274;
  assign T274 = divValidReceived_2 & T244;
  assign T275 = T277 | T276;
  assign T276 = divValidReceived_1 & T251;
  assign T277 = divValidReceived_0 & T258;
  assign T278 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T279 = 10'h3/* 3*/ == T280;
  assign T280 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T281 = ! T282;
  assign T282 = GS_step1PipeValidMove && T283;
  assign T283 = T284 == 10'h3/* 3*/;
  assign T284 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T285 = T286 || divValidReceived_3;
  assign T286 = divPort_rep_valid && T287;
  assign T287 = divPort_rep_tag == 10'h3/* 3*/;
  assign T288 = GS_step1PRegPostOff_valid_2 && GS_step1AllOffloadsValid_2;
  assign T289 = GS_step1PRegPostOff_valid_1 && GS_step1AllOffloadsValid_1;
  assign T290 = GS_step1PRegPostOff_valid_0 && GS_step1AllOffloadsValid_0;
  assign T291 = GS_step2PRegPreOff_ready || T292;
  assign T292 = ! GS_step2PRegPreOff_valid;
  assign T293 = T291 && T121;
  assign T294 = T119 ? 1'h0/* 0*/ : T295;
  assign T295 = T293 ? T296 : GS_step2PRegPreOff_valid;
  assign T296 = T298 | T297;
  assign T297 = GS_step1PRegPostOff_valid_3 & T134;
  assign T298 = T300 | T299;
  assign T299 = GS_step1PRegPostOff_valid_2 & T142;
  assign T300 = T302 | T301;
  assign T301 = GS_step1PRegPostOff_valid_1 & T168;
  assign T302 = GS_step1PRegPostOff_valid_0 & T192;
  assign T303 = T13 ? 1'h0/* 0*/ : T304;
  assign T304 = T97 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_3;
  assign T305 = ! GS_step2PRegPostOff_valid_2;
  assign T306 = T308 || T307;
  assign T307 = GS_step2PipeValidMove && T22;
  assign T308 = T101 && T309;
  assign T309 = T99[2'h2/* 2*/];
  assign T310 = T307 ? 1'h0/* 0*/ : T311;
  assign T311 = T308 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_2;
  assign T312 = ! GS_step2PRegPostOff_valid_1;
  assign T313 = T315 || T314;
  assign T314 = GS_step2PipeValidMove && T48;
  assign T315 = T101 && T316;
  assign T316 = T99[1'h1/* 1*/];
  assign T317 = T314 ? 1'h0/* 0*/ : T318;
  assign T318 = T315 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_1;
  assign T319 = ! GS_step2PRegPostOff_valid_0;
  assign T320 = T322 || T321;
  assign T321 = GS_step2PipeValidMove && T72;
  assign T322 = T101 && T323;
  assign T323 = T99[1'h0/* 0*/];
  assign T324 = T321 ? 1'h0/* 0*/ : T325;
  assign T325 = T322 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_0;
  assign T326 = T343 && T327;
  assign T327 = ! T328;
  assign T328 = T338 | T329;
  assign T329 = mulValidReceived_3 & T98;
  assign T330 = T334 && T331;
  assign T331 = mulValidReceived_3 || T332;
  assign T332 = mulPort_rep_valid && T333;
  assign T333 = mulPort_rep_tag == 10'h3/* 3*/;
  assign T334 = ! T335;
  assign T335 = GS_step2PipeValidMove && T336;
  assign T336 = T337 == 10'h3/* 3*/;
  assign T337 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T338 = T340 | T339;
  assign T339 = mulValidReceived_2 & T309;
  assign T340 = T342 | T341;
  assign T341 = mulValidReceived_1 & T316;
  assign T342 = mulValidReceived_0 & T323;
  assign T343 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T344 = 10'h3/* 3*/ == T345;
  assign T345 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T346 = ! T347;
  assign T347 = GS_step2PipeValidMove && T348;
  assign T348 = T349 == 10'h3/* 3*/;
  assign T349 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T350 = T351 || mulValidReceived_3;
  assign T351 = mulPort_rep_valid && T352;
  assign T352 = mulPort_rep_tag == 10'h3/* 3*/;
  assign T353 = GS_step2PRegPostOff_valid_2 && GS_step2AllOffloadsValid_2;
  assign T354 = GS_step2PRegPostOff_valid_1 && GS_step2AllOffloadsValid_1;
  assign T355 = GS_step2PRegPostOff_valid_0 && GS_step2AllOffloadsValid_0;
  assign T356 = outputReg_ready || T357;
  assign T357 = ! outputReg_valid;
  assign T358 = T0 || T359;
  assign T359 = T356 && T360;
  assign T360 = ! T1;
  assign T361 = T359 ? 1'h0/* 0*/ : T362;
  assign T362 = T0 ? T363 : outputReg_valid;
  assign T363 = T365 | T364;
  assign T364 = GS_step2PRegPostOff_valid_3 & T14;
  assign T365 = T367 | T366;
  assign T366 = GS_step2PRegPostOff_valid_2 & T22;
  assign T367 = T369 | T368;
  assign T368 = GS_step2PRegPostOff_valid_1 & T48;
  assign T369 = GS_step2PRegPostOff_valid_0 & T72;
  assign T371 = T0 ? T372 : outputReg_tag;
  assign T372 = T398 | T373;
  assign T373 = GS_step2PRegPostOff_tag_3 & T374;
  assign T374 = {4'ha/* 10*/{T14}};
  assign T376 = T97 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_3;
  assign T378 = T293 ? T379 : GS_step2PRegPreOff_tag;
  assign T379 = T384 | T380;
  assign T380 = GS_step1PRegPostOff_tag_3 & T381;
  assign T381 = {4'ha/* 10*/{T134}};
  assign T383 = T218 ? io_in_tag : GS_step1PRegPostOff_tag_3;
  assign T384 = T389 | T385;
  assign T385 = GS_step1PRegPostOff_tag_2 & T386;
  assign T386 = {4'ha/* 10*/{T142}};
  assign T388 = T243 ? io_in_tag : GS_step1PRegPostOff_tag_2;
  assign T389 = T394 | T390;
  assign T390 = GS_step1PRegPostOff_tag_1 & T391;
  assign T391 = {4'ha/* 10*/{T168}};
  assign T393 = T250 ? io_in_tag : GS_step1PRegPostOff_tag_1;
  assign T394 = GS_step1PRegPostOff_tag_0 & T395;
  assign T395 = {4'ha/* 10*/{T192}};
  assign T397 = T257 ? io_in_tag : GS_step1PRegPostOff_tag_0;
  assign T398 = T403 | T399;
  assign T399 = GS_step2PRegPostOff_tag_2 & T400;
  assign T400 = {4'ha/* 10*/{T22}};
  assign T402 = T308 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_2;
  assign T403 = T408 | T404;
  assign T404 = GS_step2PRegPostOff_tag_1 & T405;
  assign T405 = {4'ha/* 10*/{T48}};
  assign T407 = T315 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_1;
  assign T408 = GS_step2PRegPostOff_tag_0 & T409;
  assign T409 = {4'ha/* 10*/{T72}};
  assign T411 = T322 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_0;
  assign io_out_valid = outputReg_valid;
  assign io_in_ready = T412;
  assign T412 = GS_step1PRegPostOff_ready && GS_step1AllOffloadsReady;
  RREncode_3 GS_step1RThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T254 ),
       .io_valid_1( T247 ),
       .io_valid_2( T240 ),
       .io_valid_3( T131 ),
       .io_chosen( GS_step1RThreadEncoder_io_chosen ),
       .io_ready( GS_step1PipeReadyMove ));
  RREncode_4 GS_step1VThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T290 ),
       .io_valid_1( T289 ),
       .io_valid_2( T288 ),
       .io_valid_3( T122 ),
       .io_chosen( GS_step1VThreadEncoder_io_chosen ),
       .io_ready( GS_step1PipeValidMove ));
  RREncode_5 GS_step2RThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T319 ),
       .io_valid_1( T312 ),
       .io_valid_2( T305 ),
       .io_valid_3( T11 ),
       .io_chosen( GS_step2RThreadEncoder_io_chosen ),
       .io_ready( GS_step2PipeReadyMove ));
  RREncode_6 GS_step2VThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T355 ),
       .io_valid_1( T354 ),
       .io_valid_2( T353 ),
       .io_valid_3( T2 ),
       .io_chosen( GS_step2VThreadEncoder_io_chosen ),
       .io_ready( GS_step2PipeValidMove ));

  always @(posedge clk) begin
    if(reset) begin
      outputReg_tag <= T370;
    end else if(T0) begin
      outputReg_tag <= T371;
    end
    mulPortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T5;
    if(reset) begin
      GS_step2PRegPostOff_valid_3 <= 1'h0/* 0*/;
    end else if(T12) begin
      GS_step2PRegPostOff_valid_3 <= T303;
    end
    mulPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T25;
    mulValidReceived_2 <= reset ? 1'h0/* 0*/ : T35;
    mulPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T51;
    mulValidReceived_1 <= reset ? 1'h0/* 0*/ : T61;
    mulPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T75;
    mulValidReceived_0 <= reset ? 1'h0/* 0*/ : T85;
    mulPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T106;
    mulReadyReceived <= reset ? 1'h0/* 0*/ : T114;
    if(reset) begin
      GS_step2PRegPreOff_valid <= 1'h0/* 0*/;
    end else if(T118) begin
      GS_step2PRegPreOff_valid <= T294;
    end
    divPortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T125;
    if(reset) begin
      GS_step1PRegPostOff_valid_3 <= 1'h0/* 0*/;
    end else if(T132) begin
      GS_step1PRegPostOff_valid_3 <= T238;
    end
    divPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T145;
    divValidReceived_2 <= reset ? 1'h0/* 0*/ : T155;
    divPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T171;
    divValidReceived_1 <= reset ? 1'h0/* 0*/ : T181;
    divPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T195;
    divValidReceived_0 <= reset ? 1'h0/* 0*/ : T205;
    divPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T227;
    divReadyReceived <= reset ? 1'h0/* 0*/ : T235;
    if(reset) begin
      GS_step1PRegPostOff_valid_2 <= 1'h0/* 0*/;
    end else if(T241) begin
      GS_step1PRegPostOff_valid_2 <= T245;
    end
    if(reset) begin
      GS_step1PRegPostOff_valid_1 <= 1'h0/* 0*/;
    end else if(T248) begin
      GS_step1PRegPostOff_valid_1 <= T252;
    end
    if(reset) begin
      GS_step1PRegPostOff_valid_0 <= 1'h0/* 0*/;
    end else if(T255) begin
      GS_step1PRegPostOff_valid_0 <= T259;
    end
    divValidReceived_3 <= reset ? 1'h0/* 0*/ : T265;
    if(reset) begin
      GS_step2PRegPostOff_valid_2 <= 1'h0/* 0*/;
    end else if(T306) begin
      GS_step2PRegPostOff_valid_2 <= T310;
    end
    if(reset) begin
      GS_step2PRegPostOff_valid_1 <= 1'h0/* 0*/;
    end else if(T313) begin
      GS_step2PRegPostOff_valid_1 <= T317;
    end
    if(reset) begin
      GS_step2PRegPostOff_valid_0 <= 1'h0/* 0*/;
    end else if(T320) begin
      GS_step2PRegPostOff_valid_0 <= T324;
    end
    mulValidReceived_3 <= reset ? 1'h0/* 0*/ : T330;
    if(reset) begin
      outputReg_valid <= 1'h0/* 0*/;
    end else if(T358) begin
      outputReg_valid <= T361;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_3 <= T375;
    end else if(T97) begin
      GS_step2PRegPostOff_tag_3 <= T376;
    end
    if(reset) begin
      GS_step2PRegPreOff_tag <= T377;
    end else if(T293) begin
      GS_step2PRegPreOff_tag <= T378;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_3 <= T382;
    end else if(T218) begin
      GS_step1PRegPostOff_tag_3 <= T383;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_2 <= T387;
    end else if(T243) begin
      GS_step1PRegPostOff_tag_2 <= T388;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_1 <= T392;
    end else if(T250) begin
      GS_step1PRegPostOff_tag_1 <= T393;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_0 <= T396;
    end else if(T257) begin
      GS_step1PRegPostOff_tag_0 <= T397;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_2 <= T401;
    end else if(T308) begin
      GS_step2PRegPostOff_tag_2 <= T402;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_1 <= T406;
    end else if(T315) begin
      GS_step2PRegPostOff_tag_1 <= T407;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_0 <= T410;
    end else if(T322) begin
      GS_step2PRegPostOff_tag_0 <= T411;
    end
  end
endmodule

module gPipe(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_div_req_ready,
    output mainOff_div_req_valid,
    output[63:0] mainOff_div_req_bits_in1,
    output[63:0] mainOff_div_req_bits_in2,
    output[9:0] mainOff_div_req_tag,
    output mainOff_div_rep_ready,
    input  mainOff_div_rep_valid,
    input [63:0] mainOff_div_rep_bits_out,
    input [9:0] mainOff_div_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul_rep_ready;
  wire[9:0] mainComp_mainOff_mul_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_div_rep_ready;
  wire[9:0] mainComp_mainOff_div_req_tag;
  wire mainComp_mainOff_div_req_valid;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_div_rep_ready = mainComp_mainOff_div_rep_ready;
  assign mainOff_div_req_tag = mainComp_mainOff_div_req_tag;
  assign mainOff_div_req_valid = mainComp_mainOff_div_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  rankCalculator mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_damping( io_in_bits_damping ),
       .io_in_bits_rank(  ),
       .io_in_bits_fanoutDegree(  ),
       .io_in_tag( io_in_tag ),
       .outputReg_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mul_req_ready( offComp_io_in_ready ),
       .mainOff_mul_req_valid( mainComp_mainOff_mul_req_valid ),
       .mainOff_mul_req_bits_in1( mainComp_mainOff_mul_req_bits_in1 ),
       .mainOff_mul_req_bits_in2( mainComp_mainOff_mul_req_bits_in2 ),
       .mainOff_mul_req_tag( mainComp_mainOff_mul_req_tag ),
       .mainOff_mul_rep_ready( mainComp_mainOff_mul_rep_ready ),
       .mainOff_mul_rep_valid( offComp_io_out_valid ),
       .mainOff_mul_rep_bits_out(  ),
       .mainOff_mul_rep_tag( offComp_io_out_tag ),
       .mainOff_div_req_ready( mainOff_div_req_ready ),
       .mainOff_div_req_valid( mainComp_mainOff_div_req_valid ),
       .mainOff_div_req_bits_in1(  ),
       .mainOff_div_req_bits_in2(  ),
       .mainOff_div_req_tag( mainComp_mainOff_div_req_tag ),
       .mainOff_div_rep_ready( mainComp_mainOff_div_rep_ready ),
       .mainOff_div_rep_valid( mainOff_div_rep_valid ),
       .mainOff_div_rep_bits_out( mainOff_div_rep_bits_out ),
       .mainOff_div_rep_tag( mainOff_div_rep_tag ));
  FUSynWrapper offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul_req_tag ),
       .io_out_ready( mainComp_mainOff_mul_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_1 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_ddiv_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_div_rep_ready;
  wire[9:0] mainComp_mainOff_div_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_div_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_div_req_bits_in1;
  wire[63:0] mainComp_mainOff_div_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_damping( io_in_bits_damping ),
       .io_in_bits_rank( io_in_bits_rank ),
       .io_in_bits_fanoutDegree( io_in_bits_fanoutDegree ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_div_req_ready( offComp_io_in_ready ),
       .mainOff_div_req_valid( mainComp_mainOff_div_req_valid ),
       .mainOff_div_req_bits_in1( mainComp_mainOff_div_req_bits_in1 ),
       .mainOff_div_req_bits_in2( mainComp_mainOff_div_req_bits_in2 ),
       .mainOff_div_req_tag( mainComp_mainOff_div_req_tag ),
       .mainOff_div_rep_ready( mainComp_mainOff_div_rep_ready ),
       .mainOff_div_rep_valid( offComp_io_out_valid ),
       .mainOff_div_rep_bits_out(  ),
       .mainOff_div_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_div_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_div_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_div_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_div_req_tag ),
       .io_out_ready( mainComp_mainOff_div_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  pcIn0_valid,
    input  pcIn0_bits_request,
    input [15:0] pcIn0_bits_moduleId,
    input [7:0] pcIn0_bits_portId,
    input [19:0] pcIn0_bits_pcValue,
    input [3:0] pcIn0_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag);

  wire mainComp_mainOff_mem_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_rankCalc_rep_ready;
  wire mainComp_mainOff_rankCalc_req_valid;
  wire[9:0] mainComp_mainOff_rankCalc_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_out_bits_done;
  wire[31:0] mainComp_io_out_bits_pageId;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire offComp_io_in_ready;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_rankCalc_req_bits_damping;
  wire[31:0] mainComp_mainOff_rankCalc_req_bits_fanoutDegree;
  wire[63:0] mainComp_mainOff_rankCalc_req_bits_rank;

  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_done = mainComp_io_out_bits_done;
  assign io_out_bits_pageId = mainComp_io_out_bits_pageId;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateGenerator mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_done( mainComp_io_out_bits_done ),
       .io_out_bits_pageId( mainComp_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_rankCalc_req_ready( offComp_io_in_ready ),
       .mainOff_rankCalc_req_valid( mainComp_mainOff_rankCalc_req_valid ),
       .mainOff_rankCalc_req_bits_damping( mainComp_mainOff_rankCalc_req_bits_damping ),
       .mainOff_rankCalc_req_bits_rank( mainComp_mainOff_rankCalc_req_bits_rank ),
       .mainOff_rankCalc_req_bits_fanoutDegree( mainComp_mainOff_rankCalc_req_bits_fanoutDegree ),
       .mainOff_rankCalc_req_tag( mainComp_mainOff_rankCalc_req_tag ),
       .mainOff_rankCalc_rep_ready( mainComp_mainOff_rankCalc_rep_ready ),
       .mainOff_rankCalc_rep_valid( offComp_io_out_valid ),
       .mainOff_rankCalc_rep_bits_out(  ),
       .mainOff_rankCalc_rep_tag( offComp_io_out_tag ));
  gOffloadedComponent_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_rankCalc_req_valid ),
       .io_in_bits_damping( mainComp_mainOff_rankCalc_req_bits_damping ),
       .io_in_bits_rank( mainComp_mainOff_rankCalc_req_bits_rank ),
       .io_in_bits_fanoutDegree( mainComp_mainOff_rankCalc_req_bits_fanoutDegree ),
       .io_in_tag( mainComp_mainOff_rankCalc_req_tag ),
       .io_out_ready( mainComp_mainOff_rankCalc_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_7(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_8(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_9(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateGenerator_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_rankCalc_req_ready,
    output mainOff_rankCalc_req_valid,
    output[63:0] mainOff_rankCalc_req_bits_damping,
    output[63:0] mainOff_rankCalc_req_bits_rank,
    output[31:0] mainOff_rankCalc_req_bits_fanoutDegree,
    output[9:0] mainOff_rankCalc_req_tag,
    output mainOff_rankCalc_rep_ready,
    input  mainOff_rankCalc_rep_valid,
    input [63:0] mainOff_rankCalc_rep_bits_out,
    input [9:0] mainOff_rankCalc_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_1;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[4:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_1;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] rankCalcPortHadValidRequest_1;
  wire T12;
  wire T13;
  wire T14;
  wire rankCalcPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[4:0] T24;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_1;
  wire T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire AllOffloadsReady;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg[0:0] rankCalcPortHadReadyRequest;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg[0:0] rankCalc_ready_received;
  wire T46;
  wire T47;
  wire rankCalcPort_req_ready;
  wire rankCalcPort_rep_ready;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire memPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[7:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  reg[0:0] mem_valid_received_1;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[9:0] T75;
  wire[9:0] memPort_rep_tag;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T76;
  wire[165:0] T77;
  wire[165:0] T78;
  wire[3:0] T79;
  wire[165:0] T80;
  wire[165:0] T81;
  wire[3:0] T82;
  wire[165:0] T83;
  wire[165:0] T84;
  wire[165:0] T85;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T86;
  wire[57:0] T87;
  wire[57:0] T88;
  wire[33:0] T89;
  wire[31:0] T90;
  wire[31:0] T91;
  wire[31:0] T92;
  reg[31:0] linkId_1;
  wire T93;
  wire T94;
  wire T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire T102;
  reg[7:0] State_0;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[7:0] T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[7:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[7:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[7:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[31:0] page_fanoutDegree;
  wire[31:0] T132;
  wire[127:0] memRep1_data;
  wire[127:0] T133;
  wire[127:0] memPortReplyValue;
  wire[127:0] T134;
  wire[127:0] T135;
  wire[127:0] T136;
  wire[127:0] T137;
  reg[127:0] memPortReplyStorage_1_data;
  wire T138;
  wire T139;
  wire[1:0] T140;
  wire[1024:0] T141;
  wire memPort_rep_valid;
  wire[127:0] T142;
  wire[127:0] memPort_rep_bits_data;
  wire[127:0] T143;
  wire[127:0] T144;
  reg[127:0] memPortReplyStorage_0_data;
  wire T145;
  wire T146;
  wire[127:0] T147;
  wire[127:0] T148;
  wire T149;
  wire T150;
  wire[9:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[31:0] T157;
  wire[31:0] T158;
  wire[31:0] T159;
  wire[31:0] T160;
  wire[31:0] T161;
  reg[31:0] inputReg_1_length;
  wire T162;
  wire T163;
  wire[1:0] T164;
  wire[4:0] T165;
  wire T166;
  wire T167;
  wire[31:0] T168;
  wire[31:0] T169;
  wire[31:0] T170;
  reg[31:0] inputReg_0_length;
  wire T171;
  wire T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T176;
  reg[31:0] inputReg_1_startPageId;
  wire[31:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  reg[31:0] inputReg_0_startPageId;
  wire[31:0] T180;
  wire[31:0] T181;
  wire[31:0] T182;
  wire[31:0] T183;
  reg[31:0] pageId_1;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire[31:0] T189;
  wire[31:0] T190;
  wire T191;
  wire T192;
  wire[31:0] T193;
  wire[31:0] T194;
  wire[31:0] T195;
  reg[31:0] fanoutDegree_1;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[31:0] T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire[31:0] T206;
  wire[31:0] T207;
  reg[31:0] fanoutDegree_0;
  wire T208;
  wire T209;
  wire T210;
  wire[31:0] T211;
  wire[31:0] T212;
  wire[31:0] T213;
  wire[31:0] T214;
  wire[31:0] T215;
  reg[31:0] linkIndex_1;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire[31:0] T221;
  wire[31:0] T222;
  wire[31:0] T223;
  wire[31:0] T224;
  wire[31:0] T225;
  reg[31:0] linkIndex_0;
  wire T226;
  wire T227;
  wire[31:0] T228;
  wire[31:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[7:0] T235;
  wire T236;
  wire[31:0] T237;
  wire[31:0] T238;
  wire[31:0] T239;
  wire[31:0] T240;
  wire[31:0] T241;
  wire[31:0] T242;
  wire[31:0] T243;
  reg[31:0] pageId_0;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[7:0] T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  reg[0:0] inputReg_1_done;
  wire T273;
  wire T274;
  reg[0:0] inputReg_0_done;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  reg[0:0] outputReg_1_done;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  reg[0:0] outputReg_0_done;
  wire T293;
  wire T294;
  wire T295;
  wire[31:0] T296;
  wire[31:0] T297;
  wire[31:0] T298;
  reg[31:0] outputReg_1_pageId;
  wire T299;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[31:0] T305;
  reg[31:0] outPageId_1;
  wire T306;
  wire[127:0] T307;
  wire[127:0] T308;
  wire[127:0] T309;
  wire[127:0] T310;
  wire[127:0] T311;
  reg[127:0] memRep_1_data;
  wire T312;
  wire T313;
  wire T314;
  wire[127:0] T315;
  wire[127:0] T316;
  wire[127:0] T317;
  wire[127:0] T318;
  wire[127:0] T319;
  reg[127:0] memRep_0_data;
  wire T320;
  wire T321;
  wire T322;
  wire[127:0] T323;
  wire[127:0] T324;
  wire[127:0] T325;
  wire[31:0] T326;
  wire[31:0] T327;
  reg[31:0] outPageId_0;
  wire[127:0] T328;
  wire[127:0] T329;
  wire[31:0] T330;
  wire[31:0] T331;
  reg[31:0] outputReg_0_pageId;
  wire T332;
  wire[31:0] T333;
  wire[31:0] T334;
  wire T335;
  wire T336;
  wire T337;
  wire[7:0] T338;
  wire[7:0] T339;
  wire[7:0] T340;
  wire[7:0] T341;
  wire[7:0] T342;
  wire[7:0] T343;
  wire[7:0] T344;
  wire[7:0] T345;
  wire[7:0] T346;
  wire[7:0] T347;
  wire[7:0] T348;
  wire[7:0] T349;
  wire[7:0] T350;
  wire[7:0] T351;
  wire[7:0] T352;
  wire[7:0] T353;
  reg[7:0] EmitReturnState_1;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire[7:0] T360;
  wire[7:0] T361;
  wire[7:0] T362;
  wire[7:0] T363;
  wire[7:0] T364;
  wire[7:0] T365;
  wire[7:0] T366;
  wire[7:0] T367;
  wire[7:0] T368;
  wire[7:0] T369;
  reg[7:0] EmitReturnState_0;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[7:0] T378;
  wire[7:0] T379;
  wire[7:0] T380;
  wire[7:0] T381;
  wire[7:0] T382;
  wire[7:0] T383;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[7:0] T386;
  wire[7:0] T387;
  wire[7:0] T388;
  wire[7:0] T389;
  wire T390;
  wire T391;
  wire[127:0] T392;
  wire[127:0] T393;
  wire[127:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  reg[31:0] linkId_0;
  wire[127:0] T397;
  wire[127:0] T398;
  wire T399;
  wire T400;
  wire[7:0] T401;
  wire T402;
  wire[127:0] T403;
  wire T404;
  wire T405;
  wire[31:0] T406;
  wire[165:0] T407;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T408;
  wire[34:0] T409;
  wire[34:0] T410;
  wire[31:0] T411;
  wire[31:0] T412;
  wire[31:0] T413;
  wire[31:0] T414;
  wire[31:0] T415;
  wire[34:0] T416;
  wire T417;
  wire T418;
  wire[7:0] T419;
  wire T420;
  wire[127:0] T421;
  wire T422;
  wire T423;
  wire[31:0] T424;
  wire[165:0] T425;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T426;
  wire[55:0] T427;
  wire[55:0] T428;
  wire[34:0] T429;
  wire T430;
  wire T431;
  wire[7:0] T432;
  wire T433;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T434;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T435;
  wire memPort_req_bits_cached;
  wire T436;
  wire memPort_req_bits_rw;
  wire T437;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T438;
  wire T439;
  wire T440;
  wire[4:0] T441;
  wire T442;
  reg[0:0] mem_valid_received_0;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire[9:0] T447;
  wire T448;
  wire T449;
  wire[4:0] T450;
  wire T451;
  wire T452;
  reg[0:0] memPortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] mem_ready_received;
  wire T457;
  wire T458;
  wire memPort_req_ready;
  wire T459;
  wire T460;
  reg[0:0] subStateTh_0;
  wire T461;
  wire T462;
  wire T463;
  wire[1:0] T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire[1:0] T471;
  wire T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  reg[0:0] rankCalc_valid_received_1;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[9:0] T484;
  wire[9:0] rankCalcPort_rep_tag;
  wire[9:0] rankCalcPort_req_tag;
  wire[9:0] T485;
  wire rankCalcPort_rep_valid;
  wire T486;
  wire T487;
  wire[4:0] T488;
  wire T489;
  reg[0:0] rankCalc_valid_received_0;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[9:0] T494;
  wire T495;
  wire T496;
  wire[4:0] T497;
  wire T498;
  wire T499;
  wire[4:0] T500;
  wire T501;
  wire T502;
  wire[4:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[9:0] T507;
  wire T508;
  wire T509;
  reg[0:0] memPortHadValidRequest_1;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire[4:0] T514;
  wire T515;
  wire T516;
  wire[4:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[9:0] T521;
  wire T522;
  wire T523;
  wire AllOffloadsValid_0;
  wire T524;
  wire T525;
  wire T526;
  reg[0:0] rankCalcPortHadValidRequest_0;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire[4:0] T531;
  wire T532;
  wire T533;
  wire[4:0] T534;
  wire T535;
  wire T536;
  wire T537;
  wire[9:0] T538;
  wire T539;
  wire T540;
  reg[0:0] memPortHadValidRequest_0;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire[4:0] T545;
  wire T546;
  wire T547;
  wire[4:0] T548;
  wire T549;
  wire T550;
  wire T551;
  wire[9:0] T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire[7:0] T571;
  wire[7:0] T572;
  wire[7:0] T573;
  wire[7:0] T574;
  wire[7:0] T575;
  wire[7:0] T576;
  wire[7:0] T577;
  wire[7:0] T578;
  wire[7:0] T579;
  wire[7:0] T580;
  wire[7:0] T581;
  wire[7:0] T582;
  wire[7:0] T583;
  wire[7:0] T584;
  wire[7:0] T585;
  wire[7:0] T586;
  wire[7:0] T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[9:0] T597;
  wire[9:0] T598;
  wire[9:0] T599;
  reg[9:0] inputTag_1;
  wire[9:0] T600;
  wire[9:0] T601;
  wire[9:0] T602;
  reg[9:0] inputTag_0;
  wire[9:0] T603;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T1 = T592 && T2;
  assign T2 = State_1 == 8'h0/* 0*/;
  assign T3 = T555 || T4;
  assign T4 = T105 && T5;
  assign T5 = T6[1'h1/* 1*/];
  assign T6 = T7[1'h1/* 1*/:1'h0/* 0*/];
  assign T7 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T522 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T9;
  assign T9 = T508 && T10;
  assign T10 = T504 || T11;
  assign T11 = ! rankCalcPortHadValidRequest_1;
  assign T12 = T501 && T13;
  assign T13 = rankCalcPortHadValidRequest_1 || T14;
  assign T14 = T499 && rankCalcPort_req_valid;
  assign rankCalcPort_req_valid = T15;
  assign T15 = T476 && T16;
  assign T16 = T475 && T17;
  assign T17 = T19 == T18;
  assign T18 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T19 = T473 | T20;
  assign T20 = State_1 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23[1'h1/* 1*/];
  assign T23 = T24[1'h1/* 1*/:1'h0/* 0*/];
  assign T24 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_1 == 1'h0/* 0*/;
  assign T26 = T30 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_1;
  assign T28 = T29 == vThreadEncoder_io_chosen;
  assign T29 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T30 = T32 && T31;
  assign T31 = State_1 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_1 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = T36 == rThreadEncoder_io_chosen;
  assign T36 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign AllOffloadsReady = T37;
  assign T37 = T49 && T38;
  assign T38 = T45 || T39;
  assign T39 = T41 && T40;
  assign T40 = ! rankCalcPort_req_valid;
  assign T41 = ! rankCalcPortHadReadyRequest;
  assign T42 = T44 && T43;
  assign T43 = rankCalcPortHadReadyRequest || rankCalcPort_req_valid;
  assign T44 = ! AllOffloadsReady;
  assign T45 = rankCalcPort_req_ready || rankCalc_ready_received;
  assign T46 = T48 && T47;
  assign T47 = rankCalc_ready_received || rankCalcPort_req_ready;
  assign rankCalcPort_req_ready = mainOff_rankCalc_req_ready;
  assign mainOff_rankCalc_rep_ready = rankCalcPort_rep_ready;
  assign rankCalcPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_rankCalc_req_valid = rankCalcPort_req_valid;
  assign T48 = ! AllOffloadsReady;
  assign T49 = T456 || T50;
  assign T50 = T452 && T51;
  assign T51 = ! memPort_req_valid;
  assign memPort_req_valid = T52;
  assign T52 = T67 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T19 == T56;
  assign T56 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T19 == T61;
  assign T61 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T63 = T66 && T64;
  assign T64 = T19 == T65;
  assign T65 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T66 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T67 = T451 && T68;
  assign T68 = ! T69;
  assign T69 = T442 | T70;
  assign T70 = mem_valid_received_1 & T22;
  assign T71 = T439 && T72;
  assign T72 = mem_valid_received_1 || T73;
  assign T73 = memPort_rep_valid && T74;
  assign T74 = memPort_rep_tag == T75;
  assign T75 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T76;
  assign T76 = T77[8'ha5/* 165*/:8'h86/* 134*/];
  assign T77 = T430 ? T425 : T78;
  assign T78 = {T424, T423, T422, T421, T79};
  assign T79 = T80[2'h3/* 3*/:1'h0/* 0*/];
  assign T80 = T417 ? T407 : T81;
  assign T81 = {T406, T405, T404, T403, T82};
  assign T82 = T83[2'h3/* 3*/:1'h0/* 0*/];
  assign T83 = T399 ? T85 : T84;
  assign T84 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T85 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h4/* 4*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T86;
  assign T86 = T87[5'h1f/* 31*/:1'h0/* 0*/];
  assign T87 = 58'h4000000/* 67108864*/ + T88;
  assign T88 = {24'h0/* 0*/, T89};
  assign T89 = T90 << 32'h2/* 2*/;
  assign T90 = T395 | T91;
  assign T91 = linkId_1 & T92;
  assign T92 = {6'h20/* 32*/{T22}};
  assign T93 = T94 && T5;
  assign T94 = T391 && T95;
  assign T95 = T97 == T96;
  assign T96 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T97 = T100 | T98;
  assign T98 = State_1 & T99;
  assign T99 = {4'h8/* 8*/{T5}};
  assign T100 = State_0 & T101;
  assign T101 = {4'h8/* 8*/{T102}};
  assign T102 = T6[1'h0/* 0*/];
  assign T103 = T109 || T104;
  assign T104 = T105 && T102;
  assign T105 = T108 && T106;
  assign T106 = T97 == T107;
  assign T107 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T108 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T109 = T115 || T110;
  assign T110 = T111 && T102;
  assign T111 = T114 && T112;
  assign T112 = T97 == T113;
  assign T113 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T114 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T115 = T121 || T116;
  assign T116 = T117 && T102;
  assign T117 = T120 && T118;
  assign T118 = T97 == T119;
  assign T119 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T120 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T121 = T127 || T122;
  assign T122 = T123 && T102;
  assign T123 = T126 && T124;
  assign T124 = T97 == T125;
  assign T125 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T126 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T127 = T152 || T128;
  assign T128 = T129 && T102;
  assign T129 = T94 && T130;
  assign T130 = ! T131;
  assign T131 = page_fanoutDegree == 32'h0/* 0*/;
  assign page_fanoutDegree = T132;
  assign T132 = memRep1_data[5'h1f/* 31*/:1'h0/* 0*/];
  assign memRep1_data = T133;
  assign T133 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T149 ? T148 : T134;
  assign T134 = {T135};
  assign T135 = T143 | T136;
  assign T136 = memPortReplyStorage_1_data & T137;
  assign T137 = {8'h80/* 128*/{T5}};
  assign T138 = memPort_rep_valid && T139;
  assign T139 = T140[1'h1/* 1*/];
  assign T140 = T141[1'h1/* 1*/:1'h0/* 0*/];
  assign T141 = 2'h1/* 1*/ << memPort_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T142 = T138 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign T143 = memPortReplyStorage_0_data & T144;
  assign T144 = {8'h80/* 128*/{T102}};
  assign T145 = memPort_rep_valid && T146;
  assign T146 = T140[1'h0/* 0*/];
  assign T147 = T145 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T148 = {memPort_rep_bits_data};
  assign T149 = memPort_rep_valid && T150;
  assign T150 = T151 == memPort_rep_tag;
  assign T151 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = T252 || T153;
  assign T153 = T154 && T102;
  assign T154 = T251 && T155;
  assign T155 = ! T156;
  assign T156 = T181 == T157;
  assign T157 = T158 - 32'h1/* 1*/;
  assign T158 = T174 + T159;
  assign T159 = T169 | T160;
  assign T160 = inputReg_1_length & T161;
  assign T161 = {6'h20/* 32*/{T5}};
  assign T162 = T166 && T163;
  assign T163 = T164[1'h1/* 1*/];
  assign T164 = T165[1'h1/* 1*/:1'h0/* 0*/];
  assign T165 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T166 = T167 && io_in_valid;
  assign T167 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T168 = T162 ? io_in_bits_length : inputReg_1_length;
  assign T169 = inputReg_0_length & T170;
  assign T170 = {6'h20/* 32*/{T102}};
  assign T171 = T166 && T172;
  assign T172 = T164[1'h0/* 0*/];
  assign T173 = T171 ? io_in_bits_length : inputReg_0_length;
  assign T174 = T178 | T175;
  assign T175 = inputReg_1_startPageId & T176;
  assign T176 = {6'h20/* 32*/{T5}};
  assign T177 = T162 ? io_in_bits_startPageId : inputReg_1_startPageId;
  assign T178 = inputReg_0_startPageId & T179;
  assign T179 = {6'h20/* 32*/{T102}};
  assign T180 = T171 ? io_in_bits_startPageId : inputReg_0_startPageId;
  assign T181 = T242 | T182;
  assign T182 = pageId_1 & T183;
  assign T183 = {6'h20/* 32*/{T5}};
  assign T184 = T230 || T185;
  assign T185 = T186 && T5;
  assign T186 = T191 && T187;
  assign T187 = ! T188;
  assign T188 = T181 == T189;
  assign T189 = T190 - 32'h1/* 1*/;
  assign T190 = T174 + T159;
  assign T191 = T111 && T192;
  assign T192 = T213 == T193;
  assign T193 = T206 | T194;
  assign T194 = fanoutDegree_1 & T195;
  assign T195 = {6'h20/* 32*/{T5}};
  assign T196 = T201 || T197;
  assign T197 = T198 && T5;
  assign T198 = T94 && T199;
  assign T199 = ! T200;
  assign T200 = page_fanoutDegree <= 32'h20/* 32*/;
  assign T201 = T202 && T5;
  assign T202 = T94 && T200;
  assign T203 = T197 ? T205 : T204;
  assign T204 = T201 ? page_fanoutDegree : fanoutDegree_1;
  assign T205 = page_fanoutDegree & 32'h1f/* 31*/;
  assign T206 = fanoutDegree_0 & T207;
  assign T207 = {6'h20/* 32*/{T102}};
  assign T208 = T210 || T209;
  assign T209 = T198 && T102;
  assign T210 = T202 && T102;
  assign T211 = T209 ? T205 : T212;
  assign T212 = T210 ? page_fanoutDegree : fanoutDegree_0;
  assign T213 = T224 | T214;
  assign T214 = linkIndex_1 & T215;
  assign T215 = {6'h20/* 32*/{T5}};
  assign T216 = T220 || T217;
  assign T217 = T218 && T5;
  assign T218 = T111 && T219;
  assign T219 = ! T192;
  assign T220 = T123 && T5;
  assign T221 = T217 ? T223 : T222;
  assign T222 = T220 ? 32'h0/* 0*/ : linkIndex_1;
  assign T223 = T213 + 32'h1/* 1*/;
  assign T224 = linkIndex_0 & T225;
  assign T225 = {6'h20/* 32*/{T102}};
  assign T226 = T122 || T227;
  assign T227 = T218 && T102;
  assign T228 = T227 ? T223 : T229;
  assign T229 = T122 ? 32'h0/* 0*/ : linkIndex_0;
  assign T230 = T232 || T231;
  assign T231 = T154 && T5;
  assign T232 = T233 && T5;
  assign T233 = T236 && T234;
  assign T234 = T97 == T235;
  assign T235 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T236 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T237 = T185 ? T241 : T238;
  assign T238 = T231 ? T240 : T239;
  assign T239 = T232 ? T174 : pageId_1;
  assign T240 = T181 + 32'h1/* 1*/;
  assign T241 = T181 + 32'h1/* 1*/;
  assign T242 = pageId_0 & T243;
  assign T243 = {6'h20/* 32*/{T102}};
  assign T244 = T246 || T245;
  assign T245 = T186 && T102;
  assign T246 = T247 || T153;
  assign T247 = T233 && T102;
  assign T248 = T245 ? T241 : T249;
  assign T249 = T153 ? T240 : T250;
  assign T250 = T247 ? T174 : pageId_0;
  assign T251 = T94 && T131;
  assign T252 = T255 || T253;
  assign T253 = T254 && T102;
  assign T254 = T251 && T156;
  assign T255 = T261 || T256;
  assign T256 = T257 && T102;
  assign T257 = T260 && T258;
  assign T258 = T97 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T261 = T267 || T262;
  assign T262 = T263 && T102;
  assign T263 = T266 && T264;
  assign T264 = T97 == T265;
  assign T265 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T266 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T267 = T276 || T268;
  assign T268 = T269 && T102;
  assign T269 = T233 && T270;
  assign T270 = ! T271;
  assign T271 = T274 | T272;
  assign T272 = inputReg_1_done & T5;
  assign T273 = T162 ? io_in_bits_done : inputReg_1_done;
  assign T274 = inputReg_0_done & T102;
  assign T275 = T171 ? io_in_bits_done : inputReg_0_done;
  assign T276 = T279 || T277;
  assign T277 = T278 && T102;
  assign T278 = T233 && T271;
  assign T279 = T171 || T280;
  assign T280 = T282 && T281;
  assign T281 = T23[1'h0/* 0*/];
  assign T282 = T335 && io_out_ready;
  assign io_out_valid = T283;
  assign T283 = T285 && T284;
  assign T284 = T19 == 8'hff/* 255*/;
  assign T285 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_bits_done = T286;
  assign T286 = T292 | T287;
  assign T287 = outputReg_1_done & T22;
  assign T288 = T289 || T4;
  assign T289 = T263 && T5;
  assign T290 = T4 ? T271 : T291;
  assign T291 = T289 ? 1'h0/* 0*/ : outputReg_1_done;
  assign T292 = outputReg_0_done & T281;
  assign T293 = T262 || T104;
  assign T294 = T104 ? T271 : T295;
  assign T295 = T262 ? 1'h0/* 0*/ : outputReg_0_done;
  assign io_out_bits_pageId = T296;
  assign T296 = T330 | T297;
  assign T297 = outputReg_1_pageId & T298;
  assign T298 = {6'h20/* 32*/{T22}};
  assign T299 = T289 || T300;
  assign T300 = T111 && T5;
  assign T301 = T300 ? T303 : T302;
  assign T302 = T289 ? T181 : outputReg_1_pageId;
  assign T303 = T326 | T304;
  assign T304 = outPageId_1 & T305;
  assign T305 = {6'h20/* 32*/{T5}};
  assign T306 = T117 && T5;
  assign T307 = T306 ? T309 : T308;
  assign T308 = {96'h0/* 0*/, outPageId_1};
  assign T309 = T318 | T310;
  assign T310 = memRep_1_data & T311;
  assign T311 = {8'h80/* 128*/{T5}};
  assign T312 = T313 || T306;
  assign T313 = T314 || T93;
  assign T314 = T257 && T5;
  assign T315 = T306 ? T133 : T316;
  assign T316 = T93 ? memRep1_data : T317;
  assign T317 = T314 ? T133 : memRep_1_data;
  assign T318 = memRep_0_data & T319;
  assign T319 = {8'h80/* 128*/{T102}};
  assign T320 = T321 || T116;
  assign T321 = T256 || T322;
  assign T322 = T94 && T102;
  assign T323 = T116 ? T133 : T324;
  assign T324 = T322 ? memRep1_data : T325;
  assign T325 = T256 ? T133 : memRep_0_data;
  assign T326 = outPageId_0 & T327;
  assign T327 = {6'h20/* 32*/{T102}};
  assign T328 = T116 ? T309 : T329;
  assign T329 = {96'h0/* 0*/, outPageId_0};
  assign T330 = outputReg_0_pageId & T331;
  assign T331 = {6'h20/* 32*/{T281}};
  assign T332 = T262 || T110;
  assign T333 = T110 ? T303 : T334;
  assign T334 = T262 ? T181 : outputReg_0_pageId;
  assign T335 = T337 && T336;
  assign T336 = T19 == 8'hff/* 255*/;
  assign T337 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T338 = T390 ? 8'hff/* 255*/ : T339;
  assign T339 = T116 ? T389 : T340;
  assign T340 = T122 ? T388 : T341;
  assign T341 = T128 ? T387 : T342;
  assign T342 = T153 ? T386 : T343;
  assign T343 = T253 ? 8'h0/* 0*/ : T344;
  assign T344 = T256 ? T385 : T345;
  assign T345 = T262 ? 8'hff/* 255*/ : T346;
  assign T346 = T268 ? T384 : T347;
  assign T347 = T277 ? T383 : T348;
  assign T348 = T280 ? T351 : T349;
  assign T349 = T171 ? T350 : State_0;
  assign T350 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T351 = T368 | T352;
  assign T352 = EmitReturnState_1 & T353;
  assign T353 = {4'h8/* 8*/{T22}};
  assign T354 = T355 || T4;
  assign T355 = T356 || T217;
  assign T356 = T357 || T185;
  assign T357 = T289 || T358;
  assign T358 = T359 && T5;
  assign T359 = T191 && T188;
  assign T360 = T4 ? 8'h0/* 0*/ : T361;
  assign T361 = T217 ? T367 : T362;
  assign T362 = T185 ? T366 : T363;
  assign T363 = T358 ? 8'h0/* 0*/ : T364;
  assign T364 = T289 ? T365 : EmitReturnState_1;
  assign T365 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T366 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T367 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T368 = EmitReturnState_0 & T369;
  assign T369 = {4'h8/* 8*/{T281}};
  assign T370 = T371 || T104;
  assign T371 = T372 || T227;
  assign T372 = T373 || T245;
  assign T373 = T262 || T374;
  assign T374 = T359 && T102;
  assign T375 = T104 ? 8'h0/* 0*/ : T376;
  assign T376 = T227 ? T382 : T377;
  assign T377 = T245 ? T381 : T378;
  assign T378 = T374 ? 8'h0/* 0*/ : T379;
  assign T379 = T262 ? T380 : EmitReturnState_0;
  assign T380 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T381 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T382 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T383 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T384 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T385 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T386 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T387 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T388 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T389 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T390 = T110 || T104;
  assign T391 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T392 = T93 ? T394 : T393;
  assign T393 = {96'h0/* 0*/, linkId_1};
  assign T394 = memRep1_data >> 32'h20/* 32*/;
  assign T395 = linkId_0 & T396;
  assign T396 = {6'h20/* 32*/{T281}};
  assign T397 = T322 ? T394 : T398;
  assign T398 = {96'h0/* 0*/, linkId_0};
  assign T399 = T402 && T400;
  assign T400 = T19 == T401;
  assign T401 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T402 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T403 = T83[8'h83/* 131*/:3'h4/* 4*/];
  assign T404 = T83[8'h84/* 132*/];
  assign T405 = T83[8'h85/* 133*/];
  assign T406 = T83[8'ha5/* 165*/:8'h86/* 134*/];
  assign T407 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h8/* 8*/;
  assign memReq2_cached = 1'h0/* 0*/;
  assign memReq2_rw = 1'h0/* 0*/;
  assign memReq2_addr = T408;
  assign T408 = T409[5'h1f/* 31*/:1'h0/* 0*/];
  assign T409 = T416 + T410;
  assign T410 = T411 << 32'h3/* 3*/;
  assign T411 = T414 | T412;
  assign T412 = pageId_1 & T413;
  assign T413 = {6'h20/* 32*/{T22}};
  assign T414 = pageId_0 & T415;
  assign T415 = {6'h20/* 32*/{T281}};
  assign T416 = {3'h0/* 0*/, 32'h0/* 0*/};
  assign T417 = T420 && T418;
  assign T418 = T19 == T419;
  assign T419 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T420 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T421 = T80[8'h83/* 131*/:3'h4/* 4*/];
  assign T422 = T80[8'h84/* 132*/];
  assign T423 = T80[8'h85/* 133*/];
  assign T424 = T80[8'ha5/* 165*/:8'h86/* 134*/];
  assign T425 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h8/* 8*/;
  assign memReq1_cached = 1'h0/* 0*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T426;
  assign T426 = T427[5'h1f/* 31*/:1'h0/* 0*/];
  assign T427 = 56'h1000000/* 16777216*/ + T428;
  assign T428 = {21'h0/* 0*/, T429};
  assign T429 = T411 << 32'h3/* 3*/;
  assign T430 = T433 && T431;
  assign T431 = T19 == T432;
  assign T432 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T433 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_valid = memPort_req_valid;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T434;
  assign T434 = T77[2'h3/* 3*/:1'h0/* 0*/];
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T435;
  assign T435 = T77[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T436;
  assign T436 = T77[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T437;
  assign T437 = T77[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T438;
  assign T438 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T439 = ! T440;
  assign T440 = T441 == 5'h1/* 1*/;
  assign T441 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T442 = mem_valid_received_0 & T281;
  assign T443 = T448 && T444;
  assign T444 = mem_valid_received_0 || T445;
  assign T445 = memPort_rep_valid && T446;
  assign T446 = memPort_rep_tag == T447;
  assign T447 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T448 = ! T449;
  assign T449 = T450 == 5'h0/* 0*/;
  assign T450 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T451 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T452 = ! memPortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = memPortHadReadyRequest || memPort_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = memPort_req_ready || mem_ready_received;
  assign T457 = T459 && T458;
  assign T458 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = subStateTh_0 == 1'h0/* 0*/;
  assign T461 = T465 ? 1'h1/* 1*/ : T462;
  assign T462 = T463 ? 1'h0/* 0*/ : subStateTh_0;
  assign T463 = T464 == vThreadEncoder_io_chosen;
  assign T464 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T465 = T467 && T466;
  assign T466 = State_0 != 8'hff/* 255*/;
  assign T467 = T469 && T468;
  assign T468 = State_0 != 8'h0/* 0*/;
  assign T469 = AllOffloadsReady && T470;
  assign T470 = T471 == rThreadEncoder_io_chosen;
  assign T471 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T472 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T473 = State_0 & T474;
  assign T474 = {4'h8/* 8*/{T281}};
  assign T475 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T476 = T498 && T477;
  assign T477 = ! T478;
  assign T478 = T489 | T479;
  assign T479 = rankCalc_valid_received_1 & T22;
  assign T480 = T486 && T481;
  assign T481 = rankCalc_valid_received_1 || T482;
  assign T482 = rankCalcPort_rep_valid && T483;
  assign T483 = rankCalcPort_rep_tag == T484;
  assign T484 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign rankCalcPort_rep_tag = mainOff_rankCalc_rep_tag;
  assign mainOff_rankCalc_req_tag = rankCalcPort_req_tag;
  assign rankCalcPort_req_tag = T485;
  assign T485 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign rankCalcPort_rep_valid = mainOff_rankCalc_rep_valid;
  assign T486 = ! T487;
  assign T487 = T488 == 5'h1/* 1*/;
  assign T488 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T489 = rankCalc_valid_received_0 & T281;
  assign T490 = T495 && T491;
  assign T491 = rankCalc_valid_received_0 || T492;
  assign T492 = rankCalcPort_rep_valid && T493;
  assign T493 = rankCalcPort_rep_tag == T494;
  assign T494 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T495 = ! T496;
  assign T496 = T497 == 5'h0/* 0*/;
  assign T497 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T498 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T499 = 5'h1/* 1*/ == T500;
  assign T500 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T501 = ! T502;
  assign T502 = T503 == 5'h1/* 1*/;
  assign T503 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T504 = T505 || rankCalc_valid_received_1;
  assign T505 = rankCalcPort_rep_valid && T506;
  assign T506 = rankCalcPort_rep_tag == T507;
  assign T507 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T508 = T518 || T509;
  assign T509 = ! memPortHadValidRequest_1;
  assign T510 = T515 && T511;
  assign T511 = memPortHadValidRequest_1 || T512;
  assign T512 = T513 && memPort_req_valid;
  assign T513 = 5'h1/* 1*/ == T514;
  assign T514 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T515 = ! T516;
  assign T516 = T517 == 5'h1/* 1*/;
  assign T517 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T518 = T519 || mem_valid_received_1;
  assign T519 = memPort_rep_valid && T520;
  assign T520 = memPort_rep_tag == T521;
  assign T521 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T522 = subStateTh_1 == 1'h1/* 1*/;
  assign T523 = T553 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T524;
  assign T524 = T539 && T525;
  assign T525 = T535 || T526;
  assign T526 = ! rankCalcPortHadValidRequest_0;
  assign T527 = T532 && T528;
  assign T528 = rankCalcPortHadValidRequest_0 || T529;
  assign T529 = T530 && rankCalcPort_req_valid;
  assign T530 = 5'h0/* 0*/ == T531;
  assign T531 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T532 = ! T533;
  assign T533 = T534 == 5'h0/* 0*/;
  assign T534 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T535 = T536 || rankCalc_valid_received_0;
  assign T536 = rankCalcPort_rep_valid && T537;
  assign T537 = rankCalcPort_rep_tag == T538;
  assign T538 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T539 = T549 || T540;
  assign T540 = ! memPortHadValidRequest_0;
  assign T541 = T546 && T542;
  assign T542 = memPortHadValidRequest_0 || T543;
  assign T543 = T544 && memPort_req_valid;
  assign T544 = 5'h0/* 0*/ == T545;
  assign T545 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T546 = ! T547;
  assign T547 = T548 == 5'h0/* 0*/;
  assign T548 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T549 = T550 || mem_valid_received_0;
  assign T550 = memPort_rep_valid && T551;
  assign T551 = memPort_rep_tag == T552;
  assign T552 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T553 = subStateTh_0 == 1'h1/* 1*/;
  assign T554 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T555 = T556 || T300;
  assign T556 = T557 || T306;
  assign T557 = T558 || T220;
  assign T558 = T560 || T559;
  assign T559 = T129 && T5;
  assign T560 = T561 || T231;
  assign T561 = T563 || T562;
  assign T562 = T254 && T5;
  assign T563 = T564 || T314;
  assign T564 = T565 || T289;
  assign T565 = T567 || T566;
  assign T566 = T269 && T5;
  assign T567 = T569 || T568;
  assign T568 = T278 && T5;
  assign T569 = T162 || T570;
  assign T570 = T282 && T22;
  assign T571 = T591 ? 8'hff/* 255*/ : T572;
  assign T572 = T306 ? T590 : T573;
  assign T573 = T220 ? T589 : T574;
  assign T574 = T559 ? T588 : T575;
  assign T575 = T231 ? T587 : T576;
  assign T576 = T562 ? 8'h0/* 0*/ : T577;
  assign T577 = T314 ? T586 : T578;
  assign T578 = T289 ? 8'hff/* 255*/ : T579;
  assign T579 = T566 ? T585 : T580;
  assign T580 = T568 ? T584 : T581;
  assign T581 = T570 ? T351 : T582;
  assign T582 = T162 ? T583 : State_1;
  assign T583 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T584 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T585 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T586 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T587 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T588 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T589 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T590 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T591 = T300 || T4;
  assign T592 = subStateTh_1 == 1'h0/* 0*/;
  assign T593 = T595 && T594;
  assign T594 = State_0 == 8'h0/* 0*/;
  assign T595 = subStateTh_0 == 1'h0/* 0*/;
  assign T596 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_tag = T597;
  assign T597 = T601 | T598;
  assign T598 = inputTag_1 & T599;
  assign T599 = {4'ha/* 10*/{T22}};
  assign T600 = T162 ? io_in_tag : inputTag_1;
  assign T601 = inputTag_0 & T602;
  assign T602 = {4'ha/* 10*/{T281}};
  assign T603 = T171 ? io_in_tag : inputTag_0;
  RREncode_7 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T460 ),
       .io_valid_1( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T472 ));
  RREncode_8 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T523 ),
       .io_valid_1( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T554 ));
  RREncode_9 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T593 ),
       .io_valid_1( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T596 ));

  always @(posedge clk) begin
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_1 <= T571;
    end
    rankCalcPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T26;
    rankCalcPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T42;
    rankCalc_ready_received <= reset ? 1'h0/* 0*/ : T46;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T71;
    if(T93) begin
      linkId_1 <= T392;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T103) begin
      State_0 <= T338;
    end
    if(T138) begin
      memPortReplyStorage_1_data <= T142;
    end
    if(T145) begin
      memPortReplyStorage_0_data <= T147;
    end
    if(T162) begin
      inputReg_1_length <= T168;
    end
    if(T171) begin
      inputReg_0_length <= T173;
    end
    if(T162) begin
      inputReg_1_startPageId <= T177;
    end
    if(T171) begin
      inputReg_0_startPageId <= T180;
    end
    if(T184) begin
      pageId_1 <= T237;
    end
    if(T196) begin
      fanoutDegree_1 <= T203;
    end
    if(T208) begin
      fanoutDegree_0 <= T211;
    end
    if(T216) begin
      linkIndex_1 <= T221;
    end
    if(T226) begin
      linkIndex_0 <= T228;
    end
    if(T244) begin
      pageId_0 <= T248;
    end
    if(T162) begin
      inputReg_1_done <= T273;
    end
    if(T171) begin
      inputReg_0_done <= T275;
    end
    if(T288) begin
      outputReg_1_done <= T290;
    end
    if(T293) begin
      outputReg_0_done <= T294;
    end
    if(T299) begin
      outputReg_1_pageId <= T301;
    end
    if(T306) begin
      outPageId_1 <= T307;
    end
    if(T312) begin
      memRep_1_data <= T315;
    end
    if(T320) begin
      memRep_0_data <= T323;
    end
    if(T116) begin
      outPageId_0 <= T328;
    end
    if(T332) begin
      outputReg_0_pageId <= T333;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T354) begin
      EmitReturnState_1 <= T360;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T370) begin
      EmitReturnState_0 <= T375;
    end
    if(T322) begin
      linkId_0 <= T397;
    end
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T443;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T457;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T461;
    rankCalc_valid_received_1 <= reset ? 1'h0/* 0*/ : T480;
    rankCalc_valid_received_0 <= reset ? 1'h0/* 0*/ : T490;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T510;
    rankCalcPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T527;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T541;
    if(T162) begin
      inputTag_1 <= T600;
    end
    if(T171) begin
      inputTag_0 <= T603;
    end
  end
endmodule

module RREncode_10(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_11(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_12(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module RREncode_13(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    output[2:0] io_chosen,
    input  io_ready);

  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  reg[1:0] last_grant;
  wire T13;
  wire outValid;
  wire T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;

  assign io_chosen = choose;
  assign choose = T22 ? T21 : T0;
  assign T0 = T19 ? T18 : T1;
  assign T1 = T11 ? T10 : T2;
  assign T2 = io_valid_0 ? T9 : T3;
  assign T3 = io_valid_1 ? T8 : T4;
  assign T4 = io_valid_2 ? T7 : T5;
  assign T5 = io_valid_3 ? T6 : 3'h4/* 4*/;
  assign T6 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T7 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T8 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T9 = {2'h0/* 0*/, 1'h0/* 0*/};
  assign T10 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T11 = io_valid_3 && T12;
  assign T12 = 2'h3/* 3*/ > last_grant;
  assign T13 = outValid && io_ready;
  assign outValid = T14 || io_valid_3;
  assign T14 = T15 || io_valid_2;
  assign T15 = io_valid_0 || io_valid_1;
  assign T16 = T13 ? choose : T17;
  assign T17 = {1'h0/* 0*/, last_grant};
  assign T18 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T19 = io_valid_2 && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {2'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_valid_1 && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T13) begin
      last_grant <= T16;
    end
  end
endmodule

module rankCalculator_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  outputReg_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mul_req_ready,
    output mainOff_mul_req_valid,
    output[63:0] mainOff_mul_req_bits_in1,
    output[63:0] mainOff_mul_req_bits_in2,
    output[9:0] mainOff_mul_req_tag,
    output mainOff_mul_rep_ready,
    input  mainOff_mul_rep_valid,
    input [63:0] mainOff_mul_rep_bits_out,
    input [9:0] mainOff_mul_rep_tag,
    input  mainOff_div_req_ready,
    output mainOff_div_req_valid,
    output[63:0] mainOff_div_req_bits_in1,
    output[63:0] mainOff_div_req_bits_in2,
    output[9:0] mainOff_div_req_tag,
    output mainOff_div_rep_ready,
    input  mainOff_div_rep_valid,
    input [63:0] mainOff_div_rep_bits_out,
    input [9:0] mainOff_div_rep_tag);

  wire T0;
  wire GS_step1AllOffloadsReady;
  wire T1;
  wire T2;
  wire T3;
  wire divPort_req_valid;
  wire T4;
  wire T5;
  wire T6;
  wire[2:0] GS_step1RThreadEncoder_io_chosen;
  wire T7;
  reg[0:0] GS_step1PRegPostOff_valid_3;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[10:0] T12;
  wire[2:0] GS_step1VThreadEncoder_io_chosen;
  wire T13;
  wire GS_step1AllOffloadsValid_3;
  wire T14;
  wire T15;
  reg[0:0] divPortHadValidRequest_3;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[9:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[9:0] T24;
  wire GS_step1PipeValidMove;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire GS_step1AllOffloadsValid_2;
  wire T31;
  wire T32;
  reg[0:0] divPortHadValidRequest_2;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[9:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[9:0] T41;
  wire T42;
  reg[0:0] divValidReceived_2;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[9:0] divPort_rep_tag;
  wire divPort_rep_ready;
  wire[9:0] divPort_req_tag;
  wire[9:0] T47;
  wire divPort_rep_valid;
  wire T48;
  wire T49;
  wire T50;
  wire[9:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire GS_step1AllOffloadsValid_1;
  wire T57;
  wire T58;
  reg[0:0] divPortHadValidRequest_1;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[9:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire[9:0] T67;
  wire T68;
  reg[0:0] divValidReceived_1;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[9:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire GS_step1AllOffloadsValid_0;
  wire T81;
  wire T82;
  reg[0:0] divPortHadValidRequest_0;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[9:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[9:0] T91;
  wire T92;
  reg[0:0] divValidReceived_0;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[9:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire GS_step2PRegPreOff_ready;
  wire T104;
  wire GS_step2AllOffloadsReady;
  wire T105;
  wire T106;
  wire T107;
  wire mulPort_req_valid;
  wire T108;
  wire T109;
  wire T110;
  wire[2:0] GS_step2RThreadEncoder_io_chosen;
  wire T111;
  reg[0:0] GS_step2PRegPostOff_valid_3;
  wire T112;
  wire T113;
  wire T114;
  wire[3:0] T115;
  wire[10:0] T116;
  wire[2:0] GS_step2VThreadEncoder_io_chosen;
  wire T117;
  wire GS_step2AllOffloadsValid_3;
  wire T118;
  wire T119;
  reg[0:0] mulPortHadValidRequest_3;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire[9:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[9:0] T128;
  wire GS_step2PipeValidMove;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire GS_step2AllOffloadsValid_2;
  wire T135;
  wire T136;
  reg[0:0] mulPortHadValidRequest_2;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[9:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[9:0] T145;
  wire T146;
  reg[0:0] mulValidReceived_2;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire[9:0] mulPort_rep_tag;
  wire mulPort_rep_ready;
  wire[9:0] mulPort_req_tag;
  wire[9:0] T151;
  wire mulPort_rep_valid;
  wire T152;
  wire T153;
  wire T154;
  wire[9:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire GS_step2AllOffloadsValid_1;
  wire T161;
  wire T162;
  reg[0:0] mulPortHadValidRequest_1;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[9:0] T167;
  wire T168;
  wire T169;
  wire T170;
  wire[9:0] T171;
  wire T172;
  reg[0:0] mulValidReceived_1;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire[9:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire GS_step2AllOffloadsValid_0;
  wire T185;
  wire T186;
  reg[0:0] mulPortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[9:0] T191;
  wire T192;
  wire T193;
  wire T194;
  wire[9:0] T195;
  wire T196;
  reg[0:0] mulValidReceived_0;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[9:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  reg[0:0] mulValidReceived_3;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire[9:0] T217;
  wire T218;
  wire T219;
  wire T220;
  reg[0:0] GS_step2PRegPostOff_valid_2;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[3:0] T225;
  wire[10:0] T226;
  wire T227;
  wire T228;
  wire GS_step2PRegPostOff_ready;
  wire T229;
  reg[0:0] GS_step2PRegPreOff_valid;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  reg[0:0] GS_step1PRegPostOff_valid_2;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[3:0] T247;
  wire[10:0] T248;
  wire T249;
  wire GS_step1PRegPostOff_ready;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  reg[0:0] GS_step1PRegPostOff_valid_1;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  reg[0:0] GS_step1PRegPostOff_valid_0;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  reg[0:0] GS_step2PRegPostOff_valid_1;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  reg[0:0] GS_step2PRegPostOff_valid_0;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire GS_step2PipeReadyMove;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  reg[0:0] mulPortHadReadyRequest;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  reg[0:0] mulReadyReceived;
  wire T309;
  wire T310;
  wire mulPort_req_ready;
  wire T311;
  wire T312;
  wire T313;
  reg[0:0] divValidReceived_3;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[9:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire GS_step1PipeReadyMove;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  reg[0:0] divPortHadReadyRequest;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  reg[0:0] divReadyReceived;
  wire T352;
  wire T353;
  wire divPort_req_ready;
  wire T354;
  reg[9:0] outputReg_tag;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  reg[0:0] outputReg_valid;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire[9:0] T371;
  wire[9:0] T372;
  wire[9:0] T373;
  wire[9:0] T374;
  wire[9:0] T375;
  reg[9:0] GS_step2PRegPostOff_tag_3;
  wire[9:0] T376;
  wire[9:0] T377;
  reg[9:0] GS_step2PRegPreOff_tag;
  wire[9:0] T378;
  wire[9:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire[9:0] T382;
  reg[9:0] GS_step1PRegPostOff_tag_3;
  wire[9:0] T383;
  wire[9:0] T384;
  wire[9:0] T385;
  wire[9:0] T386;
  wire[9:0] T387;
  reg[9:0] GS_step1PRegPostOff_tag_2;
  wire[9:0] T388;
  wire[9:0] T389;
  wire[9:0] T390;
  wire[9:0] T391;
  wire[9:0] T392;
  reg[9:0] GS_step1PRegPostOff_tag_1;
  wire[9:0] T393;
  wire[9:0] T394;
  wire[9:0] T395;
  wire[9:0] T396;
  reg[9:0] GS_step1PRegPostOff_tag_0;
  wire[9:0] T397;
  wire[9:0] T398;
  wire[9:0] T399;
  wire[9:0] T400;
  wire[9:0] T401;
  reg[9:0] GS_step2PRegPostOff_tag_2;
  wire[9:0] T402;
  wire[9:0] T403;
  wire[9:0] T404;
  wire[9:0] T405;
  wire[9:0] T406;
  reg[9:0] GS_step2PRegPostOff_tag_1;
  wire[9:0] T407;
  wire[9:0] T408;
  wire[9:0] T409;
  wire[9:0] T410;
  reg[9:0] GS_step2PRegPostOff_tag_0;
  wire[9:0] T411;
  wire[9:0] T412;

  assign io_in_ready = T0;
  assign T0 = GS_step1PRegPostOff_ready && GS_step1AllOffloadsReady;
  assign GS_step1AllOffloadsReady = T1;
  assign T1 = T351 || T2;
  assign T2 = T347 && T3;
  assign T3 = ! divPort_req_valid;
  assign divPort_req_valid = T4;
  assign T4 = T337 && T5;
  assign T5 = io_in_valid && T6;
  assign T6 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T7 = ! GS_step1PRegPostOff_valid_3;
  assign T8 = T327 || T9;
  assign T9 = GS_step1PipeValidMove && T10;
  assign T10 = T11[2'h3/* 3*/];
  assign T11 = T12[2'h3/* 3*/:1'h0/* 0*/];
  assign T12 = 4'h1/* 1*/ << GS_step1VThreadEncoder_io_chosen;
  assign T13 = GS_step1PRegPostOff_valid_3 && GS_step1AllOffloadsValid_3;
  assign GS_step1AllOffloadsValid_3 = T14;
  assign T14 = T313 || T15;
  assign T15 = ! divPortHadValidRequest_3;
  assign T16 = T21 && T17;
  assign T17 = divPortHadValidRequest_3 || T18;
  assign T18 = T19 && divPort_req_valid;
  assign T19 = 10'h3/* 3*/ == T20;
  assign T20 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T21 = ! T22;
  assign T22 = GS_step1PipeValidMove && T23;
  assign T23 = T24 == 10'h3/* 3*/;
  assign T24 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign GS_step1PipeValidMove = T25;
  assign T25 = T103 && T26;
  assign T26 = T28 | T27;
  assign T27 = GS_step1AllOffloadsValid_3 & T10;
  assign T28 = T54 | T29;
  assign T29 = GS_step1AllOffloadsValid_2 & T30;
  assign T30 = T11[2'h2/* 2*/];
  assign GS_step1AllOffloadsValid_2 = T31;
  assign T31 = T42 || T32;
  assign T32 = ! divPortHadValidRequest_2;
  assign T33 = T38 && T34;
  assign T34 = divPortHadValidRequest_2 || T35;
  assign T35 = T36 && divPort_req_valid;
  assign T36 = 10'h2/* 2*/ == T37;
  assign T37 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T38 = ! T39;
  assign T39 = GS_step1PipeValidMove && T40;
  assign T40 = T41 == 10'h2/* 2*/;
  assign T41 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T42 = T52 || divValidReceived_2;
  assign T43 = T48 && T44;
  assign T44 = divValidReceived_2 || T45;
  assign T45 = divPort_rep_valid && T46;
  assign T46 = divPort_rep_tag == 10'h2/* 2*/;
  assign divPort_rep_tag = mainOff_div_rep_tag;
  assign mainOff_div_rep_ready = divPort_rep_ready;
  assign divPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_div_req_tag = divPort_req_tag;
  assign divPort_req_tag = T47;
  assign T47 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign divPort_rep_valid = mainOff_div_rep_valid;
  assign mainOff_div_req_valid = divPort_req_valid;
  assign T48 = ! T49;
  assign T49 = GS_step1PipeValidMove && T50;
  assign T50 = T51 == 10'h2/* 2*/;
  assign T51 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T52 = divPort_rep_valid && T53;
  assign T53 = divPort_rep_tag == 10'h2/* 2*/;
  assign T54 = T79 | T55;
  assign T55 = GS_step1AllOffloadsValid_1 & T56;
  assign T56 = T11[1'h1/* 1*/];
  assign GS_step1AllOffloadsValid_1 = T57;
  assign T57 = T68 || T58;
  assign T58 = ! divPortHadValidRequest_1;
  assign T59 = T64 && T60;
  assign T60 = divPortHadValidRequest_1 || T61;
  assign T61 = T62 && divPort_req_valid;
  assign T62 = 10'h1/* 1*/ == T63;
  assign T63 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T64 = ! T65;
  assign T65 = GS_step1PipeValidMove && T66;
  assign T66 = T67 == 10'h1/* 1*/;
  assign T67 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T68 = T77 || divValidReceived_1;
  assign T69 = T73 && T70;
  assign T70 = divValidReceived_1 || T71;
  assign T71 = divPort_rep_valid && T72;
  assign T72 = divPort_rep_tag == 10'h1/* 1*/;
  assign T73 = ! T74;
  assign T74 = GS_step1PipeValidMove && T75;
  assign T75 = T76 == 10'h1/* 1*/;
  assign T76 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T77 = divPort_rep_valid && T78;
  assign T78 = divPort_rep_tag == 10'h1/* 1*/;
  assign T79 = GS_step1AllOffloadsValid_0 & T80;
  assign T80 = T11[1'h0/* 0*/];
  assign GS_step1AllOffloadsValid_0 = T81;
  assign T81 = T92 || T82;
  assign T82 = ! divPortHadValidRequest_0;
  assign T83 = T88 && T84;
  assign T84 = divPortHadValidRequest_0 || T85;
  assign T85 = T86 && divPort_req_valid;
  assign T86 = 10'h0/* 0*/ == T87;
  assign T87 = {7'h0/* 0*/, GS_step1RThreadEncoder_io_chosen};
  assign T88 = ! T89;
  assign T89 = GS_step1PipeValidMove && T90;
  assign T90 = T91 == 10'h0/* 0*/;
  assign T91 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T92 = T101 || divValidReceived_0;
  assign T93 = T97 && T94;
  assign T94 = divValidReceived_0 || T95;
  assign T95 = divPort_rep_valid && T96;
  assign T96 = divPort_rep_tag == 10'h0/* 0*/;
  assign T97 = ! T98;
  assign T98 = GS_step1PipeValidMove && T99;
  assign T99 = T100 == 10'h0/* 0*/;
  assign T100 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T101 = divPort_rep_valid && T102;
  assign T102 = divPort_rep_tag == 10'h0/* 0*/;
  assign T103 = T312 && GS_step2PRegPreOff_ready;
  assign GS_step2PRegPreOff_ready = T104;
  assign T104 = GS_step2PRegPostOff_ready && GS_step2AllOffloadsReady;
  assign GS_step2AllOffloadsReady = T105;
  assign T105 = T308 || T106;
  assign T106 = T304 && T107;
  assign T107 = ! mulPort_req_valid;
  assign mulPort_req_valid = T108;
  assign T108 = T294 && T109;
  assign T109 = GS_step2PRegPreOff_valid && T110;
  assign T110 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T111 = ! GS_step2PRegPostOff_valid_3;
  assign T112 = T284 || T113;
  assign T113 = GS_step2PipeValidMove && T114;
  assign T114 = T115[2'h3/* 3*/];
  assign T115 = T116[2'h3/* 3*/:1'h0/* 0*/];
  assign T116 = 4'h1/* 1*/ << GS_step2VThreadEncoder_io_chosen;
  assign T117 = GS_step2PRegPostOff_valid_3 && GS_step2AllOffloadsValid_3;
  assign GS_step2AllOffloadsValid_3 = T118;
  assign T118 = T209 || T119;
  assign T119 = ! mulPortHadValidRequest_3;
  assign T120 = T125 && T121;
  assign T121 = mulPortHadValidRequest_3 || T122;
  assign T122 = T123 && mulPort_req_valid;
  assign T123 = 10'h3/* 3*/ == T124;
  assign T124 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T125 = ! T126;
  assign T126 = GS_step2PipeValidMove && T127;
  assign T127 = T128 == 10'h3/* 3*/;
  assign T128 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign GS_step2PipeValidMove = T129;
  assign T129 = T207 && T130;
  assign T130 = T132 | T131;
  assign T131 = GS_step2AllOffloadsValid_3 & T114;
  assign T132 = T158 | T133;
  assign T133 = GS_step2AllOffloadsValid_2 & T134;
  assign T134 = T115[2'h2/* 2*/];
  assign GS_step2AllOffloadsValid_2 = T135;
  assign T135 = T146 || T136;
  assign T136 = ! mulPortHadValidRequest_2;
  assign T137 = T142 && T138;
  assign T138 = mulPortHadValidRequest_2 || T139;
  assign T139 = T140 && mulPort_req_valid;
  assign T140 = 10'h2/* 2*/ == T141;
  assign T141 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T142 = ! T143;
  assign T143 = GS_step2PipeValidMove && T144;
  assign T144 = T145 == 10'h2/* 2*/;
  assign T145 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T146 = T156 || mulValidReceived_2;
  assign T147 = T152 && T148;
  assign T148 = mulValidReceived_2 || T149;
  assign T149 = mulPort_rep_valid && T150;
  assign T150 = mulPort_rep_tag == 10'h2/* 2*/;
  assign mulPort_rep_tag = mainOff_mul_rep_tag;
  assign mainOff_mul_rep_ready = mulPort_rep_ready;
  assign mulPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul_req_tag = mulPort_req_tag;
  assign mulPort_req_tag = T151;
  assign T151 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign mulPort_rep_valid = mainOff_mul_rep_valid;
  assign mainOff_mul_req_valid = mulPort_req_valid;
  assign T152 = ! T153;
  assign T153 = GS_step2PipeValidMove && T154;
  assign T154 = T155 == 10'h2/* 2*/;
  assign T155 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T156 = mulPort_rep_valid && T157;
  assign T157 = mulPort_rep_tag == 10'h2/* 2*/;
  assign T158 = T183 | T159;
  assign T159 = GS_step2AllOffloadsValid_1 & T160;
  assign T160 = T115[1'h1/* 1*/];
  assign GS_step2AllOffloadsValid_1 = T161;
  assign T161 = T172 || T162;
  assign T162 = ! mulPortHadValidRequest_1;
  assign T163 = T168 && T164;
  assign T164 = mulPortHadValidRequest_1 || T165;
  assign T165 = T166 && mulPort_req_valid;
  assign T166 = 10'h1/* 1*/ == T167;
  assign T167 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T168 = ! T169;
  assign T169 = GS_step2PipeValidMove && T170;
  assign T170 = T171 == 10'h1/* 1*/;
  assign T171 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T172 = T181 || mulValidReceived_1;
  assign T173 = T177 && T174;
  assign T174 = mulValidReceived_1 || T175;
  assign T175 = mulPort_rep_valid && T176;
  assign T176 = mulPort_rep_tag == 10'h1/* 1*/;
  assign T177 = ! T178;
  assign T178 = GS_step2PipeValidMove && T179;
  assign T179 = T180 == 10'h1/* 1*/;
  assign T180 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T181 = mulPort_rep_valid && T182;
  assign T182 = mulPort_rep_tag == 10'h1/* 1*/;
  assign T183 = GS_step2AllOffloadsValid_0 & T184;
  assign T184 = T115[1'h0/* 0*/];
  assign GS_step2AllOffloadsValid_0 = T185;
  assign T185 = T196 || T186;
  assign T186 = ! mulPortHadValidRequest_0;
  assign T187 = T192 && T188;
  assign T188 = mulPortHadValidRequest_0 || T189;
  assign T189 = T190 && mulPort_req_valid;
  assign T190 = 10'h0/* 0*/ == T191;
  assign T191 = {7'h0/* 0*/, GS_step2RThreadEncoder_io_chosen};
  assign T192 = ! T193;
  assign T193 = GS_step2PipeValidMove && T194;
  assign T194 = T195 == 10'h0/* 0*/;
  assign T195 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T196 = T205 || mulValidReceived_0;
  assign T197 = T201 && T198;
  assign T198 = mulValidReceived_0 || T199;
  assign T199 = mulPort_rep_valid && T200;
  assign T200 = mulPort_rep_tag == 10'h0/* 0*/;
  assign T201 = ! T202;
  assign T202 = GS_step2PipeValidMove && T203;
  assign T203 = T204 == 10'h0/* 0*/;
  assign T204 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T205 = mulPort_rep_valid && T206;
  assign T206 = mulPort_rep_tag == 10'h0/* 0*/;
  assign T207 = T208 && outputReg_ready;
  assign T208 = GS_step2VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T209 = T218 || mulValidReceived_3;
  assign T210 = T214 && T211;
  assign T211 = mulValidReceived_3 || T212;
  assign T212 = mulPort_rep_valid && T213;
  assign T213 = mulPort_rep_tag == 10'h3/* 3*/;
  assign T214 = ! T215;
  assign T215 = GS_step2PipeValidMove && T216;
  assign T216 = T217 == 10'h3/* 3*/;
  assign T217 = {7'h0/* 0*/, GS_step2VThreadEncoder_io_chosen};
  assign T218 = mulPort_rep_valid && T219;
  assign T219 = mulPort_rep_tag == 10'h3/* 3*/;
  assign T220 = GS_step2PRegPostOff_valid_2 && GS_step2AllOffloadsValid_2;
  assign T221 = T223 || T222;
  assign T222 = GS_step2PipeValidMove && T134;
  assign T223 = T227 && T224;
  assign T224 = T225[2'h2/* 2*/];
  assign T225 = T226[2'h3/* 3*/:1'h0/* 0*/];
  assign T226 = 4'h1/* 1*/ << GS_step2RThreadEncoder_io_chosen;
  assign T227 = T228 && GS_step2AllOffloadsReady;
  assign T228 = GS_step2PRegPreOff_valid && GS_step2PRegPostOff_ready;
  assign GS_step2PRegPostOff_ready = T229;
  assign T229 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T230 = T236 || T231;
  assign T231 = T234 && T232;
  assign T232 = ! T233;
  assign T233 = GS_step1VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T234 = GS_step2PRegPreOff_ready || T235;
  assign T235 = ! GS_step2PRegPreOff_valid;
  assign T236 = T234 && T233;
  assign T237 = T231 ? 1'h0/* 0*/ : T238;
  assign T238 = T236 ? T239 : GS_step2PRegPreOff_valid;
  assign T239 = T241 | T240;
  assign T240 = GS_step1PRegPostOff_valid_3 & T10;
  assign T241 = T253 | T242;
  assign T242 = GS_step1PRegPostOff_valid_2 & T30;
  assign T243 = T245 || T244;
  assign T244 = GS_step1PipeValidMove && T30;
  assign T245 = T249 && T246;
  assign T246 = T247[2'h2/* 2*/];
  assign T247 = T248[2'h3/* 3*/:1'h0/* 0*/];
  assign T248 = 4'h1/* 1*/ << GS_step1RThreadEncoder_io_chosen;
  assign T249 = GS_step1PRegPostOff_ready && GS_step1AllOffloadsReady;
  assign GS_step1PRegPostOff_ready = T250;
  assign T250 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T251 = T244 ? 1'h0/* 0*/ : T252;
  assign T252 = T245 ? io_in_valid : GS_step1PRegPostOff_valid_2;
  assign T253 = T261 | T254;
  assign T254 = GS_step1PRegPostOff_valid_1 & T56;
  assign T255 = T257 || T256;
  assign T256 = GS_step1PipeValidMove && T56;
  assign T257 = T249 && T258;
  assign T258 = T247[1'h1/* 1*/];
  assign T259 = T256 ? 1'h0/* 0*/ : T260;
  assign T260 = T257 ? io_in_valid : GS_step1PRegPostOff_valid_1;
  assign T261 = GS_step1PRegPostOff_valid_0 & T80;
  assign T262 = T264 || T263;
  assign T263 = GS_step1PipeValidMove && T80;
  assign T264 = T249 && T265;
  assign T265 = T247[1'h0/* 0*/];
  assign T266 = T263 ? 1'h0/* 0*/ : T267;
  assign T267 = T264 ? io_in_valid : GS_step1PRegPostOff_valid_0;
  assign T268 = T222 ? 1'h0/* 0*/ : T269;
  assign T269 = T223 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_2;
  assign T270 = GS_step2PRegPostOff_valid_1 && GS_step2AllOffloadsValid_1;
  assign T271 = T273 || T272;
  assign T272 = GS_step2PipeValidMove && T160;
  assign T273 = T227 && T274;
  assign T274 = T225[1'h1/* 1*/];
  assign T275 = T272 ? 1'h0/* 0*/ : T276;
  assign T276 = T273 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_1;
  assign T277 = GS_step2PRegPostOff_valid_0 && GS_step2AllOffloadsValid_0;
  assign T278 = T280 || T279;
  assign T279 = GS_step2PipeValidMove && T184;
  assign T280 = T227 && T281;
  assign T281 = T225[1'h0/* 0*/];
  assign T282 = T279 ? 1'h0/* 0*/ : T283;
  assign T283 = T280 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_0;
  assign T284 = T227 && T285;
  assign T285 = T225[2'h3/* 3*/];
  assign T286 = T113 ? 1'h0/* 0*/ : T287;
  assign T287 = T284 ? GS_step2PRegPreOff_valid : GS_step2PRegPostOff_valid_3;
  assign T288 = ! GS_step2PRegPostOff_valid_2;
  assign T289 = ! GS_step2PRegPostOff_valid_1;
  assign T290 = ! GS_step2PRegPostOff_valid_0;
  assign GS_step2PipeReadyMove = T291;
  assign T291 = T292 && GS_step2AllOffloadsReady;
  assign T292 = T293 && GS_step2PRegPostOff_ready;
  assign T293 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T294 = T303 && T295;
  assign T295 = ! T296;
  assign T296 = T298 | T297;
  assign T297 = mulValidReceived_3 & T285;
  assign T298 = T300 | T299;
  assign T299 = mulValidReceived_2 & T224;
  assign T300 = T302 | T301;
  assign T301 = mulValidReceived_1 & T274;
  assign T302 = mulValidReceived_0 & T281;
  assign T303 = GS_step2RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T304 = ! mulPortHadReadyRequest;
  assign T305 = T307 && T306;
  assign T306 = mulPortHadReadyRequest || mulPort_req_valid;
  assign T307 = ! GS_step2PipeReadyMove;
  assign T308 = mulPort_req_ready || mulReadyReceived;
  assign T309 = T311 && T310;
  assign T310 = mulReadyReceived || mulPort_req_ready;
  assign mulPort_req_ready = mainOff_mul_req_ready;
  assign T311 = ! GS_step2PipeReadyMove;
  assign T312 = GS_step1VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T313 = T322 || divValidReceived_3;
  assign T314 = T318 && T315;
  assign T315 = divValidReceived_3 || T316;
  assign T316 = divPort_rep_valid && T317;
  assign T317 = divPort_rep_tag == 10'h3/* 3*/;
  assign T318 = ! T319;
  assign T319 = GS_step1PipeValidMove && T320;
  assign T320 = T321 == 10'h3/* 3*/;
  assign T321 = {7'h0/* 0*/, GS_step1VThreadEncoder_io_chosen};
  assign T322 = divPort_rep_valid && T323;
  assign T323 = divPort_rep_tag == 10'h3/* 3*/;
  assign T324 = GS_step1PRegPostOff_valid_2 && GS_step1AllOffloadsValid_2;
  assign T325 = GS_step1PRegPostOff_valid_1 && GS_step1AllOffloadsValid_1;
  assign T326 = GS_step1PRegPostOff_valid_0 && GS_step1AllOffloadsValid_0;
  assign T327 = T249 && T328;
  assign T328 = T247[2'h3/* 3*/];
  assign T329 = T9 ? 1'h0/* 0*/ : T330;
  assign T330 = T327 ? io_in_valid : GS_step1PRegPostOff_valid_3;
  assign T331 = ! GS_step1PRegPostOff_valid_2;
  assign T332 = ! GS_step1PRegPostOff_valid_1;
  assign T333 = ! GS_step1PRegPostOff_valid_0;
  assign GS_step1PipeReadyMove = T334;
  assign T334 = T335 && GS_step1AllOffloadsReady;
  assign T335 = T336 && GS_step1PRegPostOff_ready;
  assign T336 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T337 = T346 && T338;
  assign T338 = ! T339;
  assign T339 = T341 | T340;
  assign T340 = divValidReceived_3 & T328;
  assign T341 = T343 | T342;
  assign T342 = divValidReceived_2 & T246;
  assign T343 = T345 | T344;
  assign T344 = divValidReceived_1 & T258;
  assign T345 = divValidReceived_0 & T265;
  assign T346 = GS_step1RThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T347 = ! divPortHadReadyRequest;
  assign T348 = T350 && T349;
  assign T349 = divPortHadReadyRequest || divPort_req_valid;
  assign T350 = ! GS_step1PipeReadyMove;
  assign T351 = divPort_req_ready || divReadyReceived;
  assign T352 = T354 && T353;
  assign T353 = divReadyReceived || divPort_req_ready;
  assign divPort_req_ready = mainOff_div_req_ready;
  assign T354 = ! GS_step1PipeReadyMove;
  assign io_out_tag = outputReg_tag;
  assign T355 = T357 && T356;
  assign T356 = GS_step2VThreadEncoder_io_chosen != 3'h4/* 4*/;
  assign T357 = outputReg_ready || T358;
  assign T358 = ! outputReg_valid;
  assign T359 = T355 || T360;
  assign T360 = T357 && T361;
  assign T361 = ! T356;
  assign T362 = T360 ? 1'h0/* 0*/ : T363;
  assign T363 = T355 ? T364 : outputReg_valid;
  assign T364 = T366 | T365;
  assign T365 = GS_step2PRegPostOff_valid_3 & T114;
  assign T366 = T368 | T367;
  assign T367 = GS_step2PRegPostOff_valid_2 & T134;
  assign T368 = T370 | T369;
  assign T369 = GS_step2PRegPostOff_valid_1 & T160;
  assign T370 = GS_step2PRegPostOff_valid_0 & T184;
  assign T372 = T355 ? T373 : outputReg_tag;
  assign T373 = T399 | T374;
  assign T374 = GS_step2PRegPostOff_tag_3 & T375;
  assign T375 = {4'ha/* 10*/{T114}};
  assign T377 = T284 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_3;
  assign T379 = T236 ? T380 : GS_step2PRegPreOff_tag;
  assign T380 = T385 | T381;
  assign T381 = GS_step1PRegPostOff_tag_3 & T382;
  assign T382 = {4'ha/* 10*/{T10}};
  assign T384 = T327 ? io_in_tag : GS_step1PRegPostOff_tag_3;
  assign T385 = T390 | T386;
  assign T386 = GS_step1PRegPostOff_tag_2 & T387;
  assign T387 = {4'ha/* 10*/{T30}};
  assign T389 = T245 ? io_in_tag : GS_step1PRegPostOff_tag_2;
  assign T390 = T395 | T391;
  assign T391 = GS_step1PRegPostOff_tag_1 & T392;
  assign T392 = {4'ha/* 10*/{T56}};
  assign T394 = T257 ? io_in_tag : GS_step1PRegPostOff_tag_1;
  assign T395 = GS_step1PRegPostOff_tag_0 & T396;
  assign T396 = {4'ha/* 10*/{T80}};
  assign T398 = T264 ? io_in_tag : GS_step1PRegPostOff_tag_0;
  assign T399 = T404 | T400;
  assign T400 = GS_step2PRegPostOff_tag_2 & T401;
  assign T401 = {4'ha/* 10*/{T134}};
  assign T403 = T223 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_2;
  assign T404 = T409 | T405;
  assign T405 = GS_step2PRegPostOff_tag_1 & T406;
  assign T406 = {4'ha/* 10*/{T160}};
  assign T408 = T273 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_1;
  assign T409 = GS_step2PRegPostOff_tag_0 & T410;
  assign T410 = {4'ha/* 10*/{T184}};
  assign T412 = T280 ? GS_step2PRegPreOff_tag : GS_step2PRegPostOff_tag_0;
  assign io_out_valid = outputReg_valid;
  RREncode_10 GS_step1RThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T333 ),
       .io_valid_1( T332 ),
       .io_valid_2( T331 ),
       .io_valid_3( T7 ),
       .io_chosen( GS_step1RThreadEncoder_io_chosen ),
       .io_ready( GS_step1PipeReadyMove ));
  RREncode_11 GS_step1VThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T326 ),
       .io_valid_1( T325 ),
       .io_valid_2( T324 ),
       .io_valid_3( T13 ),
       .io_chosen( GS_step1VThreadEncoder_io_chosen ),
       .io_ready( GS_step1PipeValidMove ));
  RREncode_12 GS_step2RThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T290 ),
       .io_valid_1( T289 ),
       .io_valid_2( T288 ),
       .io_valid_3( T111 ),
       .io_chosen( GS_step2RThreadEncoder_io_chosen ),
       .io_ready( GS_step2PipeReadyMove ));
  RREncode_13 GS_step2VThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T277 ),
       .io_valid_1( T270 ),
       .io_valid_2( T220 ),
       .io_valid_3( T117 ),
       .io_chosen( GS_step2VThreadEncoder_io_chosen ),
       .io_ready( GS_step2PipeValidMove ));

  always @(posedge clk) begin
    if(reset) begin
      GS_step1PRegPostOff_valid_3 <= 1'h0/* 0*/;
    end else if(T8) begin
      GS_step1PRegPostOff_valid_3 <= T329;
    end
    divPortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T16;
    divPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T33;
    divValidReceived_2 <= reset ? 1'h0/* 0*/ : T43;
    divPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T59;
    divValidReceived_1 <= reset ? 1'h0/* 0*/ : T69;
    divPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T83;
    divValidReceived_0 <= reset ? 1'h0/* 0*/ : T93;
    if(reset) begin
      GS_step2PRegPostOff_valid_3 <= 1'h0/* 0*/;
    end else if(T112) begin
      GS_step2PRegPostOff_valid_3 <= T286;
    end
    mulPortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T120;
    mulPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T137;
    mulValidReceived_2 <= reset ? 1'h0/* 0*/ : T147;
    mulPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T163;
    mulValidReceived_1 <= reset ? 1'h0/* 0*/ : T173;
    mulPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mulValidReceived_0 <= reset ? 1'h0/* 0*/ : T197;
    mulValidReceived_3 <= reset ? 1'h0/* 0*/ : T210;
    if(reset) begin
      GS_step2PRegPostOff_valid_2 <= 1'h0/* 0*/;
    end else if(T221) begin
      GS_step2PRegPostOff_valid_2 <= T268;
    end
    if(reset) begin
      GS_step2PRegPreOff_valid <= 1'h0/* 0*/;
    end else if(T230) begin
      GS_step2PRegPreOff_valid <= T237;
    end
    if(reset) begin
      GS_step1PRegPostOff_valid_2 <= 1'h0/* 0*/;
    end else if(T243) begin
      GS_step1PRegPostOff_valid_2 <= T251;
    end
    if(reset) begin
      GS_step1PRegPostOff_valid_1 <= 1'h0/* 0*/;
    end else if(T255) begin
      GS_step1PRegPostOff_valid_1 <= T259;
    end
    if(reset) begin
      GS_step1PRegPostOff_valid_0 <= 1'h0/* 0*/;
    end else if(T262) begin
      GS_step1PRegPostOff_valid_0 <= T266;
    end
    if(reset) begin
      GS_step2PRegPostOff_valid_1 <= 1'h0/* 0*/;
    end else if(T271) begin
      GS_step2PRegPostOff_valid_1 <= T275;
    end
    if(reset) begin
      GS_step2PRegPostOff_valid_0 <= 1'h0/* 0*/;
    end else if(T278) begin
      GS_step2PRegPostOff_valid_0 <= T282;
    end
    mulPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T305;
    mulReadyReceived <= reset ? 1'h0/* 0*/ : T309;
    divValidReceived_3 <= reset ? 1'h0/* 0*/ : T314;
    divPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T348;
    divReadyReceived <= reset ? 1'h0/* 0*/ : T352;
    if(reset) begin
      outputReg_tag <= T371;
    end else if(T355) begin
      outputReg_tag <= T372;
    end
    if(reset) begin
      outputReg_valid <= 1'h0/* 0*/;
    end else if(T359) begin
      outputReg_valid <= T362;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_3 <= T376;
    end else if(T284) begin
      GS_step2PRegPostOff_tag_3 <= T377;
    end
    if(reset) begin
      GS_step2PRegPreOff_tag <= T378;
    end else if(T236) begin
      GS_step2PRegPreOff_tag <= T379;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_3 <= T383;
    end else if(T327) begin
      GS_step1PRegPostOff_tag_3 <= T384;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_2 <= T388;
    end else if(T245) begin
      GS_step1PRegPostOff_tag_2 <= T389;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_1 <= T393;
    end else if(T257) begin
      GS_step1PRegPostOff_tag_1 <= T394;
    end
    if(reset) begin
      GS_step1PRegPostOff_tag_0 <= T397;
    end else if(T264) begin
      GS_step1PRegPostOff_tag_0 <= T398;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_2 <= T402;
    end else if(T223) begin
      GS_step2PRegPostOff_tag_2 <= T403;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_1 <= T407;
    end else if(T273) begin
      GS_step2PRegPostOff_tag_1 <= T408;
    end
    if(reset) begin
      GS_step2PRegPostOff_tag_0 <= T411;
    end else if(T280) begin
      GS_step2PRegPostOff_tag_0 <= T412;
    end
  end
endmodule

module gPipe_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_2 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_div_req_ready,
    output mainOff_div_req_valid,
    output[63:0] mainOff_div_req_bits_in1,
    output[63:0] mainOff_div_req_bits_in2,
    output[9:0] mainOff_div_req_tag,
    output mainOff_div_rep_ready,
    input  mainOff_div_rep_valid,
    input [63:0] mainOff_div_rep_bits_out,
    input [9:0] mainOff_div_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_div_rep_ready;
  wire[9:0] mainComp_mainOff_div_req_tag;
  wire mainComp_mainOff_div_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul_rep_ready;
  wire[9:0] mainComp_mainOff_mul_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul_req_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;
  wire[63:0] mainComp_mainOff_mul_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_div_rep_ready = mainComp_mainOff_div_rep_ready;
  assign mainOff_div_req_tag = mainComp_mainOff_div_req_tag;
  assign mainOff_div_req_valid = mainComp_mainOff_div_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  rankCalculator_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_damping( io_in_bits_damping ),
       .io_in_bits_rank(  ),
       .io_in_bits_fanoutDegree(  ),
       .io_in_tag( io_in_tag ),
       .outputReg_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mul_req_ready( offComp_io_in_ready ),
       .mainOff_mul_req_valid( mainComp_mainOff_mul_req_valid ),
       .mainOff_mul_req_bits_in1( mainComp_mainOff_mul_req_bits_in1 ),
       .mainOff_mul_req_bits_in2( mainComp_mainOff_mul_req_bits_in2 ),
       .mainOff_mul_req_tag( mainComp_mainOff_mul_req_tag ),
       .mainOff_mul_rep_ready( mainComp_mainOff_mul_rep_ready ),
       .mainOff_mul_rep_valid( offComp_io_out_valid ),
       .mainOff_mul_rep_bits_out(  ),
       .mainOff_mul_rep_tag( offComp_io_out_tag ),
       .mainOff_div_req_ready( mainOff_div_req_ready ),
       .mainOff_div_req_valid( mainComp_mainOff_div_req_valid ),
       .mainOff_div_req_bits_in1(  ),
       .mainOff_div_req_bits_in2(  ),
       .mainOff_div_req_tag( mainComp_mainOff_div_req_tag ),
       .mainOff_div_rep_ready( mainComp_mainOff_div_rep_ready ),
       .mainOff_div_rep_valid( mainOff_div_rep_valid ),
       .mainOff_div_rep_bits_out( mainOff_div_rep_bits_out ),
       .mainOff_div_rep_tag( mainOff_div_rep_tag ));
  FUSynWrapper_2 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul_req_tag ),
       .io_out_ready( mainComp_mainOff_mul_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_3 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_ddiv_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_damping,
    input [63:0] io_in_bits_rank,
    input [31:0] io_in_bits_fanoutDegree,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_div_rep_ready;
  wire[9:0] mainComp_mainOff_div_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_div_req_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;
  wire[63:0] mainComp_mainOff_div_req_bits_in1;
  wire[63:0] mainComp_mainOff_div_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_3 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_damping( io_in_bits_damping ),
       .io_in_bits_rank( io_in_bits_rank ),
       .io_in_bits_fanoutDegree( io_in_bits_fanoutDegree ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_div_req_ready( offComp_io_in_ready ),
       .mainOff_div_req_valid( mainComp_mainOff_div_req_valid ),
       .mainOff_div_req_bits_in1( mainComp_mainOff_div_req_bits_in1 ),
       .mainOff_div_req_bits_in2( mainComp_mainOff_div_req_bits_in2 ),
       .mainOff_div_req_tag( mainComp_mainOff_div_req_tag ),
       .mainOff_div_rep_ready( mainComp_mainOff_div_rep_ready ),
       .mainOff_div_rep_valid( offComp_io_out_valid ),
       .mainOff_div_rep_bits_out(  ),
       .mainOff_div_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_3 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_div_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_div_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_div_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_div_req_tag ),
       .io_out_ready( mainComp_mainOff_div_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output pcOutN_valid,
    output pcOutN_bits_request,
    output[15:0] pcOutN_bits_moduleId,
    output[7:0] pcOutN_bits_portId,
    output[19:0] pcOutN_bits_pcValue,
    output[3:0] pcOutN_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_rankCalc_rep_ready;
  wire mainComp_mainOff_rankCalc_req_valid;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire mainComp_io_out_valid;
  wire mainComp_io_out_bits_done;
  wire[31:0] mainComp_io_out_bits_pageId;
  wire mainComp_mainOff_mem_req_valid;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_rankCalc_req_tag;
  wire offComp_io_out_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_rankCalc_req_bits_damping;
  wire[31:0] mainComp_mainOff_rankCalc_req_bits_fanoutDegree;
  wire[63:0] mainComp_mainOff_rankCalc_req_bits_rank;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_done = mainComp_io_out_bits_done;
  assign io_out_bits_pageId = mainComp_io_out_bits_pageId;
  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateGenerator_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_done( mainComp_io_out_bits_done ),
       .io_out_bits_pageId( mainComp_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_rankCalc_req_ready( offComp_io_in_ready ),
       .mainOff_rankCalc_req_valid( mainComp_mainOff_rankCalc_req_valid ),
       .mainOff_rankCalc_req_bits_damping( mainComp_mainOff_rankCalc_req_bits_damping ),
       .mainOff_rankCalc_req_bits_rank( mainComp_mainOff_rankCalc_req_bits_rank ),
       .mainOff_rankCalc_req_bits_fanoutDegree( mainComp_mainOff_rankCalc_req_bits_fanoutDegree ),
       .mainOff_rankCalc_req_tag( mainComp_mainOff_rankCalc_req_tag ),
       .mainOff_rankCalc_rep_ready( mainComp_mainOff_rankCalc_rep_ready ),
       .mainOff_rankCalc_rep_valid( offComp_io_out_valid ),
       .mainOff_rankCalc_rep_bits_out(  ),
       .mainOff_rankCalc_rep_tag( offComp_io_out_tag ));
  gOffloadedComponent_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_rankCalc_req_valid ),
       .io_in_bits_damping( mainComp_mainOff_rankCalc_req_bits_damping ),
       .io_in_bits_rank( mainComp_mainOff_rankCalc_req_bits_rank ),
       .io_in_bits_fanoutDegree( mainComp_mainOff_rankCalc_req_bits_fanoutDegree ),
       .io_in_tag( mainComp_mainOff_rankCalc_req_tag ),
       .io_out_ready( mainComp_mainOff_rankCalc_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gRRDistributor(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_done,
    output[31:0] io_out_0_bits_startPageId,
    output[31:0] io_out_0_bits_length,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_done,
    output[31:0] io_out_1_bits_startPageId,
    output[31:0] io_out_1_bits_length,
    output[9:0] io_out_1_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    output io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg[0:0] last_grant;
  wire T8;
  wire T9;
  wire choose;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;

  assign io_in_ready = T0;
  assign T0 = io_out_0_ready || io_out_1_ready;
  assign io_out_1_valid = T1;
  assign T1 = T2 && io_in_valid;
  assign T2 = T15 || T3;
  assign T3 = ! T4;
  assign T4 = T5 || io_out_0_ready;
  assign T5 = T13 || T6;
  assign T6 = io_out_1_ready && T7;
  assign T7 = 1'h1/* 1*/ > last_grant;
  assign T8 = io_in_valid && io_in_ready;
  assign T9 = T8 ? choose : last_grant;
  assign choose = T11 ? 1'h1/* 1*/ : T10;
  assign T10 = io_out_0_ready ? 1'h0/* 0*/ : 1'h1/* 1*/;
  assign T11 = io_out_1_ready && T12;
  assign T12 = 1'h1/* 1*/ > last_grant;
  assign T13 = io_out_0_ready && T14;
  assign T14 = 1'h0/* 0*/ > last_grant;
  assign T15 = T17 && T16;
  assign T16 = 1'h1/* 1*/ > last_grant;
  assign T17 = ! T13;
  assign io_out_1_bits_length = io_in_bits_length;
  assign io_out_1_bits_startPageId = io_in_bits_startPageId;
  assign io_out_1_bits_done = io_in_bits_done;
  assign io_out_0_valid = T18;
  assign T18 = T19 && io_in_valid;
  assign T19 = T22 || T20;
  assign T20 = ! T21;
  assign T21 = T13 || T6;
  assign T22 = 1'h0/* 0*/ > last_grant;
  assign io_out_0_bits_done = io_in_bits_done;
  assign io_out_0_bits_length = io_in_bits_length;
  assign io_out_0_bits_startPageId = io_in_bits_startPageId;
  assign io_out_1_tag = io_in_tag;
  assign io_out_0_tag = io_in_tag;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T9;
    end
  end
endmodule

module RRDistributorComponent(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_done,
    output[31:0] io_out_0_bits_startPageId,
    output[31:0] io_out_0_bits_length,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_done,
    output[31:0] io_out_1_bits_startPageId,
    output[31:0] io_out_1_bits_length,
    output[9:0] io_out_1_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    output io_chosen);

  wire rrDist_io_in_ready;
  wire rrDist_io_out_1_valid;
  wire[31:0] rrDist_io_out_1_bits_length;
  wire[31:0] rrDist_io_out_1_bits_startPageId;
  wire rrDist_io_out_1_bits_done;
  wire rrDist_io_out_0_valid;
  wire rrDist_io_out_0_bits_done;
  wire[31:0] rrDist_io_out_0_bits_length;
  wire[31:0] rrDist_io_out_0_bits_startPageId;
  wire[9:0] rrDist_io_out_1_tag;
  wire[9:0] rrDist_io_out_0_tag;

  assign io_in_ready = rrDist_io_in_ready;
  assign io_out_1_valid = rrDist_io_out_1_valid;
  assign io_out_1_bits_length = rrDist_io_out_1_bits_length;
  assign io_out_1_bits_startPageId = rrDist_io_out_1_bits_startPageId;
  assign io_out_1_bits_done = rrDist_io_out_1_bits_done;
  assign io_out_0_valid = rrDist_io_out_0_valid;
  assign io_out_0_bits_done = rrDist_io_out_0_bits_done;
  assign io_out_0_bits_length = rrDist_io_out_0_bits_length;
  assign io_out_0_bits_startPageId = rrDist_io_out_0_bits_startPageId;
  assign io_out_1_tag = rrDist_io_out_1_tag;
  assign io_out_0_tag = rrDist_io_out_0_tag;
  gRRDistributor rrDist(.clk(clk), .reset(reset),
       .io_out_0_ready( io_out_0_ready ),
       .io_out_0_valid( rrDist_io_out_0_valid ),
       .io_out_0_bits_done( rrDist_io_out_0_bits_done ),
       .io_out_0_bits_startPageId( rrDist_io_out_0_bits_startPageId ),
       .io_out_0_bits_length( rrDist_io_out_0_bits_length ),
       .io_out_0_tag( rrDist_io_out_0_tag ),
       .io_out_1_ready( io_out_1_ready ),
       .io_out_1_valid( rrDist_io_out_1_valid ),
       .io_out_1_bits_done( rrDist_io_out_1_bits_done ),
       .io_out_1_bits_startPageId( rrDist_io_out_1_bits_startPageId ),
       .io_out_1_bits_length( rrDist_io_out_1_bits_length ),
       .io_out_1_tag( rrDist_io_out_1_tag ),
       .io_in_ready( rrDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
endmodule

module gRRArbiter(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_done,
    input [31:0] io_in_0_bits_pageId,
    input [63:0] io_in_0_bits_rankUpdate,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_done,
    input [31:0] io_in_1_bits_pageId,
    input [63:0] io_in_1_bits_rankUpdate,
    input [9:0] io_in_1_tag,
    output io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[1:0] T5;
  wire[2:0] T6;
  wire choose;
  wire T7;
  wire T8;
  wire T9;
  reg[0:0] last_grant;
  wire T10;
  wire T11;
  wire dvec_1_done;
  wire T12;
  wire T13;
  wire dvec_0_done;
  wire[31:0] T14;
  wire[31:0] T15;
  wire[31:0] T16;
  wire[31:0] dvec_1_pageId;
  wire[31:0] T17;
  wire[31:0] T18;
  wire[31:0] dvec_0_pageId;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[9:0] T35;
  wire[4:0] T36;
  wire[4:0] T37;
  wire[4:0] T38;
  wire T39;
  wire[1:0] T40;
  wire[2:0] T41;
  wire[4:0] tvec_1;
  wire[4:0] T42;
  wire[4:0] T43;
  wire[4:0] T44;
  wire T45;
  wire[4:0] tvec_0;
  wire[4:0] T46;

  assign io_in_1_ready = T0;
  assign T0 = T19 && io_out_ready;
  assign io_out_valid = T1;
  assign T1 = io_in_0_valid || io_in_1_valid;
  assign io_out_bits_done = T2;
  assign T2 = T12 | T3;
  assign T3 = dvec_1_done & T4;
  assign T4 = T5[1'h1/* 1*/];
  assign T5 = T6[1'h1/* 1*/:1'h0/* 0*/];
  assign T6 = 2'h1/* 1*/ << choose;
  assign choose = T8 ? 1'h1/* 1*/ : T7;
  assign T7 = io_in_0_valid ? 1'h0/* 0*/ : 1'h1/* 1*/;
  assign T8 = io_in_1_valid && T9;
  assign T9 = 1'h1/* 1*/ > last_grant;
  assign T10 = io_out_valid && io_out_ready;
  assign T11 = T10 ? choose : last_grant;
  assign dvec_1_done = io_in_1_bits_done;
  assign T12 = dvec_0_done & T13;
  assign T13 = T5[1'h0/* 0*/];
  assign dvec_0_done = io_in_0_bits_done;
  assign io_out_bits_pageId = T14;
  assign T14 = T17 | T15;
  assign T15 = dvec_1_pageId & T16;
  assign T16 = {6'h20/* 32*/{T4}};
  assign dvec_1_pageId = io_in_1_bits_pageId;
  assign T17 = dvec_0_pageId & T18;
  assign T18 = {6'h20/* 32*/{T13}};
  assign dvec_0_pageId = io_in_0_bits_pageId;
  assign T19 = T27 || T20;
  assign T20 = ! T21;
  assign T21 = T22 || io_in_0_valid;
  assign T22 = T25 || T23;
  assign T23 = io_in_1_valid && T24;
  assign T24 = 1'h1/* 1*/ > last_grant;
  assign T25 = io_in_0_valid && T26;
  assign T26 = 1'h0/* 0*/ > last_grant;
  assign T27 = T29 && T28;
  assign T28 = 1'h1/* 1*/ > last_grant;
  assign T29 = ! T25;
  assign io_in_0_ready = T30;
  assign T30 = T31 && io_out_ready;
  assign T31 = T34 || T32;
  assign T32 = ! T33;
  assign T33 = T25 || T23;
  assign T34 = 1'h0/* 0*/ > last_grant;
  assign io_out_tag = T35;
  assign T35 = {5'h0/* 0*/, T36};
  assign T36 = T43 | T37;
  assign T37 = tvec_1 & T38;
  assign T38 = {3'h5/* 5*/{T39}};
  assign T39 = T40[1'h1/* 1*/];
  assign T40 = T41[1'h1/* 1*/:1'h0/* 0*/];
  assign T41 = 2'h1/* 1*/ << choose;
  assign tvec_1 = T42;
  assign T42 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T43 = tvec_0 & T44;
  assign T44 = {3'h5/* 5*/{T45}};
  assign T45 = T40[1'h0/* 0*/];
  assign tvec_0 = T46;
  assign T46 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T10) begin
      last_grant <= T11;
    end
  end
endmodule

module RRAggregatorComponent(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_done,
    input [31:0] io_in_0_bits_pageId,
    input [63:0] io_in_0_bits_rankUpdate,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_done,
    input [31:0] io_in_1_bits_pageId,
    input [63:0] io_in_1_bits_rankUpdate,
    input [9:0] io_in_1_tag,
    output io_chosen);

  wire rrArb_io_in_1_ready;
  wire rrArb_io_out_valid;
  wire rrArb_io_out_bits_done;
  wire[31:0] rrArb_io_out_bits_pageId;
  wire rrArb_io_in_0_ready;
  wire[9:0] rrArb_io_out_tag;

  assign io_in_1_ready = rrArb_io_in_1_ready;
  assign io_out_valid = rrArb_io_out_valid;
  assign io_out_bits_done = rrArb_io_out_bits_done;
  assign io_out_bits_pageId = rrArb_io_out_bits_pageId;
  assign io_in_0_ready = rrArb_io_in_0_ready;
  assign io_out_tag = rrArb_io_out_tag;
  gRRArbiter rrArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( rrArb_io_out_valid ),
       .io_out_bits_done( rrArb_io_out_bits_done ),
       .io_out_bits_pageId( rrArb_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( rrArb_io_out_tag ),
       .io_in_0_ready( rrArb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_valid ),
       .io_in_0_bits_done( io_in_0_bits_done ),
       .io_in_0_bits_pageId( io_in_0_bits_pageId ),
       .io_in_0_bits_rankUpdate(  ),
       .io_in_0_tag( io_in_0_tag ),
       .io_in_1_ready( rrArb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_valid ),
       .io_in_1_bits_done( io_in_1_bits_done ),
       .io_in_1_bits_pageId( io_in_1_bits_pageId ),
       .io_in_1_bits_rankUpdate(  ),
       .io_in_1_tag( io_in_1_tag ),
       .io_chosen(  ));
endmodule

module gTaggedRRArbiter(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_addr,
    output io_out_bits_rw,
    output io_out_bits_cached,
    output[127:0] io_out_bits_data,
    output[3:0] io_out_bits_size,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_addr,
    input  io_in_0_bits_rw,
    input  io_in_0_bits_cached,
    input [127:0] io_in_0_bits_data,
    input [3:0] io_in_0_bits_size,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_addr,
    input  io_in_1_bits_rw,
    input  io_in_1_bits_cached,
    input [127:0] io_in_1_bits_data,
    input [3:0] io_in_1_bits_size,
    input [9:0] io_in_1_tag,
    output io_chosen);

  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[2:0] T5;
  wire choose;
  wire T6;
  wire[31:0] T7;
  wire[31:0] T8;
  wire[31:0] T9;
  wire[31:0] dvec_1_addr;
  wire[31:0] T10;
  wire[31:0] T11;
  wire T12;
  wire[31:0] dvec_0_addr;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg[0:0] last_grant;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] dvec_1_size;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] dvec_0_size;
  wire[127:0] T29;
  wire[127:0] T30;
  wire[127:0] T31;
  wire[127:0] dvec_1_data;
  wire[127:0] T32;
  wire[127:0] T33;
  wire[127:0] dvec_0_data;
  wire T34;
  wire T35;
  wire dvec_1_cached;
  wire T36;
  wire dvec_0_cached;
  wire T37;
  wire T38;
  wire dvec_1_rw;
  wire T39;
  wire dvec_0_rw;
  wire[9:0] T40;
  wire[6:0] T41;
  wire[6:0] T42;
  wire[6:0] T43;
  wire[4:0] T44;
  wire[4:0] T45;
  wire[4:0] T46;
  wire[4:0] tvec_1;
  wire[4:0] T47;
  wire[4:0] T48;
  wire[4:0] T49;
  wire[4:0] tvec_0;
  wire[4:0] T50;
  wire[6:0] T51;
  wire[5:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;

  assign io_out_bits_size = T0;
  assign T0 = T27 | T1;
  assign T1 = dvec_1_size & T2;
  assign T2 = {3'h4/* 4*/{T3}};
  assign T3 = T4[1'h1/* 1*/];
  assign T4 = T5[1'h1/* 1*/:1'h0/* 0*/];
  assign T5 = 2'h1/* 1*/ << choose;
  assign choose = T25 ? 1'h1/* 1*/ : T6;
  assign T6 = io_in_0_valid ? 1'h0/* 0*/ : 1'h1/* 1*/;
  assign io_out_bits_addr = T7;
  assign T7 = T10 | T8;
  assign T8 = dvec_1_addr & T9;
  assign T9 = {6'h20/* 32*/{T3}};
  assign dvec_1_addr = io_in_1_bits_addr;
  assign T10 = dvec_0_addr & T11;
  assign T11 = {6'h20/* 32*/{T12}};
  assign T12 = T4[1'h0/* 0*/];
  assign dvec_0_addr = io_in_0_bits_addr;
  assign io_out_valid = T13;
  assign T13 = io_in_0_valid || io_in_1_valid;
  assign io_in_0_ready = T14;
  assign T14 = T15 && io_out_ready;
  assign T15 = T24 || T16;
  assign T16 = ! T17;
  assign T17 = T22 || T18;
  assign T18 = io_in_1_valid && T19;
  assign T19 = 1'h1/* 1*/ > last_grant;
  assign T20 = io_out_valid && io_out_ready;
  assign T21 = T20 ? choose : last_grant;
  assign T22 = io_in_0_valid && T23;
  assign T23 = 1'h0/* 0*/ > last_grant;
  assign T24 = 1'h0/* 0*/ > last_grant;
  assign T25 = io_in_1_valid && T26;
  assign T26 = 1'h1/* 1*/ > last_grant;
  assign dvec_1_size = io_in_1_bits_size;
  assign T27 = dvec_0_size & T28;
  assign T28 = {3'h4/* 4*/{T12}};
  assign dvec_0_size = io_in_0_bits_size;
  assign io_out_bits_data = T29;
  assign T29 = T32 | T30;
  assign T30 = dvec_1_data & T31;
  assign T31 = {8'h80/* 128*/{T3}};
  assign dvec_1_data = io_in_1_bits_data;
  assign T32 = dvec_0_data & T33;
  assign T33 = {8'h80/* 128*/{T12}};
  assign dvec_0_data = io_in_0_bits_data;
  assign io_out_bits_cached = T34;
  assign T34 = T36 | T35;
  assign T35 = dvec_1_cached & T3;
  assign dvec_1_cached = io_in_1_bits_cached;
  assign T36 = dvec_0_cached & T12;
  assign dvec_0_cached = io_in_0_bits_cached;
  assign io_out_bits_rw = T37;
  assign T37 = T39 | T38;
  assign T38 = dvec_1_rw & T3;
  assign dvec_1_rw = io_in_1_bits_rw;
  assign T39 = dvec_0_rw & T12;
  assign dvec_0_rw = io_in_0_bits_rw;
  assign io_out_tag = T40;
  assign T40 = {3'h0/* 0*/, T41};
  assign T41 = T51 | T42;
  assign T42 = T43 & 7'h1f/* 31*/;
  assign T43 = {2'h0/* 0*/, T44};
  assign T44 = T48 | T45;
  assign T45 = tvec_1 & T46;
  assign T46 = {3'h5/* 5*/{T3}};
  assign tvec_1 = T47;
  assign T47 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T48 = tvec_0 & T49;
  assign T49 = {3'h5/* 5*/{T12}};
  assign tvec_0 = T50;
  assign T50 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T51 = {1'h0/* 0*/, T52};
  assign T52 = choose << 3'h5/* 5*/;
  assign io_in_1_ready = T53;
  assign T53 = T54 && io_out_ready;
  assign T54 = T58 || T55;
  assign T55 = ! T56;
  assign T56 = T57 || io_in_0_valid;
  assign T57 = T22 || T18;
  assign T58 = T60 && T59;
  assign T59 = 1'h1/* 1*/ > last_grant;
  assign T60 = ! T22;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T20) begin
      last_grant <= T21;
    end
  end
endmodule

module gTaggedDistributor(
    input  io_out_0_ready,
    output io_out_0_valid,
    output[127:0] io_out_0_bits_data,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[127:0] io_out_1_bits_data,
    output[9:0] io_out_1_tag,
    output io_in_ready,
    input  io_in_valid,
    input [127:0] io_in_bits_data,
    input [9:0] io_in_tag,
    output io_chosen);

  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T2;
  wire[9:0] T3;
  wire T4;
  wire T5;
  wire[9:0] T6;
  wire[9:0] T7;
  wire[9:0] T8;
  wire[9:0] T9;
  wire T10;
  wire T11;
  wire[9:0] T12;
  wire[9:0] T13;
  wire[9:0] T14;
  wire[9:0] T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1024:0] T21;
  wire[9:0] T22;
  wire[9:0] T23;
  wire[9:0] T24;
  wire T25;
  wire T26;

  assign io_out_1_tag = T0;
  assign T0 = io_in_tag & T1;
  assign T1 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_0_tag = T2;
  assign T2 = io_in_tag & T3;
  assign T3 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_0_valid = T4;
  assign T4 = io_in_valid && T5;
  assign T5 = T9 == T6;
  assign T6 = T8 & T7;
  assign T7 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T8 = io_in_tag >> 3'h5/* 5*/;
  assign T9 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign io_out_0_bits_data = io_in_bits_data;
  assign io_out_1_valid = T10;
  assign T10 = io_in_valid && T11;
  assign T11 = T15 == T12;
  assign T12 = T14 & T13;
  assign T13 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T14 = io_in_tag >> 3'h5/* 5*/;
  assign T15 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign io_out_1_bits_data = io_in_bits_data;
  assign io_in_ready = T16;
  assign T16 = io_in_valid && T17;
  assign T17 = T25 | T18;
  assign T18 = io_out_1_ready & T19;
  assign T19 = T20[1'h1/* 1*/];
  assign T20 = T21[1'h1/* 1*/:1'h0/* 0*/];
  assign T21 = 2'h1/* 1*/ << T22;
  assign T22 = T24 & T23;
  assign T23 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T24 = io_in_tag >> 3'h5/* 5*/;
  assign T25 = io_out_0_ready & T26;
  assign T26 = T20[1'h0/* 0*/];
endmodule

module gReplicatedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag);

  wire inputDist_io_in_ready;
  wire gOffloadedComponent_1_io_in_ready;
  wire[9:0] gTaggedDistributor_io_out_1_tag;
  wire[3:0] gTaggedRRArbiter_io_out_bits_size;
  wire gOffloadedComponent_io_off_mem_req_valid;
  wire[9:0] gTaggedDistributor_io_out_0_tag;
  wire gTaggedDistributor_io_out_0_valid;
  wire[127:0] gTaggedDistributor_io_out_0_bits_data;
  wire[31:0] gTaggedRRArbiter_io_out_bits_addr;
  wire[31:0] gOffloadedComponent_1_io_off_mem_req_bits_addr;
  wire gTaggedDistributor_io_out_1_valid;
  wire[127:0] gTaggedDistributor_io_out_1_bits_data;
  wire inputDist_io_out_1_valid;
  wire gOffloadedComponent_io_in_ready;
  wire[31:0] inputDist_io_out_1_bits_length;
  wire[31:0] inputDist_io_out_1_bits_startPageId;
  wire inputDist_io_out_1_bits_done;
  wire outputArb_io_in_1_ready;
  wire outputArb_io_out_valid;
  wire gOffloadedComponent_1_io_out_valid;
  wire gOffloadedComponent_io_out_valid;
  wire outputArb_io_out_bits_done;
  wire gOffloadedComponent_1_io_out_bits_done;
  wire gOffloadedComponent_io_out_bits_done;
  wire inputDist_io_out_0_valid;
  wire inputDist_io_out_0_bits_done;
  wire[31:0] outputArb_io_out_bits_pageId;
  wire[31:0] gOffloadedComponent_1_io_out_bits_pageId;
  wire[31:0] gOffloadedComponent_io_out_bits_pageId;
  wire[31:0] inputDist_io_out_0_bits_length;
  wire[31:0] inputDist_io_out_0_bits_startPageId;
  wire[31:0] gOffloadedComponent_io_off_mem_req_bits_addr;
  wire gTaggedRRArbiter_io_out_valid;
  wire gOffloadedComponent_1_io_off_mem_req_valid;
  wire outputArb_io_in_0_ready;
  wire gTaggedRRArbiter_io_in_0_ready;
  wire[3:0] gOffloadedComponent_1_io_off_mem_req_bits_size;
  wire[3:0] gOffloadedComponent_io_off_mem_req_bits_size;
  wire[127:0] gTaggedRRArbiter_io_out_bits_data;
  wire[127:0] gOffloadedComponent_1_io_off_mem_req_bits_data;
  wire[127:0] gOffloadedComponent_io_off_mem_req_bits_data;
  wire gTaggedRRArbiter_io_out_bits_cached;
  wire gOffloadedComponent_1_io_off_mem_req_bits_cached;
  wire gOffloadedComponent_io_off_mem_req_bits_cached;
  wire gTaggedRRArbiter_io_out_bits_rw;
  wire gOffloadedComponent_1_io_off_mem_req_bits_rw;
  wire gOffloadedComponent_io_off_mem_req_bits_rw;
  wire gTaggedDistributor_io_in_ready;
  wire gOffloadedComponent_1_io_off_mem_rep_ready;
  wire gOffloadedComponent_io_off_mem_rep_ready;
  wire[9:0] gTaggedRRArbiter_io_out_tag;
  wire[9:0] gOffloadedComponent_1_io_off_mem_req_tag;
  wire[9:0] gOffloadedComponent_io_off_mem_req_tag;
  wire gTaggedRRArbiter_io_in_1_ready;
  wire[9:0] outputArb_io_out_tag;
  wire[9:0] gOffloadedComponent_1_io_out_tag;
  wire[9:0] inputDist_io_out_1_tag;
  wire[9:0] gOffloadedComponent_io_out_tag;
  wire[9:0] inputDist_io_out_0_tag;

  assign io_in_ready = inputDist_io_in_ready;
  assign mainOff_mem_req_bits_size = gTaggedRRArbiter_io_out_bits_size;
  assign mainOff_mem_req_bits_addr = gTaggedRRArbiter_io_out_bits_addr;
  assign io_out_valid = outputArb_io_out_valid;
  assign io_out_bits_done = outputArb_io_out_bits_done;
  assign io_out_bits_pageId = outputArb_io_out_bits_pageId;
  assign mainOff_mem_req_valid = gTaggedRRArbiter_io_out_valid;
  assign mainOff_mem_req_bits_data = gTaggedRRArbiter_io_out_bits_data;
  assign mainOff_mem_req_bits_cached = gTaggedRRArbiter_io_out_bits_cached;
  assign mainOff_mem_req_bits_rw = gTaggedRRArbiter_io_out_bits_rw;
  assign mainOff_mem_rep_ready = gTaggedDistributor_io_in_ready;
  assign mainOff_mem_req_tag = gTaggedRRArbiter_io_out_tag;
  assign io_out_tag = outputArb_io_out_tag;
  gOffloadedComponent_2 gOffloadedComponent(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_io_in_ready ),
       .io_in_valid( inputDist_io_out_0_valid ),
       .io_in_bits_done( inputDist_io_out_0_bits_done ),
       .io_in_bits_startPageId( inputDist_io_out_0_bits_startPageId ),
       .io_in_bits_length( inputDist_io_out_0_bits_length ),
       .io_in_tag( inputDist_io_out_0_tag ),
       .io_out_ready( outputArb_io_in_0_ready ),
       .io_out_valid( gOffloadedComponent_io_out_valid ),
       .io_out_bits_done( gOffloadedComponent_io_out_bits_done ),
       .io_out_bits_pageId( gOffloadedComponent_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( gOffloadedComponent_io_out_tag ),
       .pcIn0_valid(  ),
       .pcIn0_bits_request(  ),
       .pcIn0_bits_moduleId(  ),
       .pcIn0_bits_portId(  ),
       .pcIn0_bits_pcValue(  ),
       .pcIn0_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_0_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_0_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_0_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_0_tag ));
  gOffloadedComponent_5 gOffloadedComponent_1(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_1_io_in_ready ),
       .io_in_valid( inputDist_io_out_1_valid ),
       .io_in_bits_done( inputDist_io_out_1_bits_done ),
       .io_in_bits_startPageId( inputDist_io_out_1_bits_startPageId ),
       .io_in_bits_length( inputDist_io_out_1_bits_length ),
       .io_in_tag( inputDist_io_out_1_tag ),
       .io_out_ready( outputArb_io_in_1_ready ),
       .io_out_valid( gOffloadedComponent_1_io_out_valid ),
       .io_out_bits_done( gOffloadedComponent_1_io_out_bits_done ),
       .io_out_bits_pageId( gOffloadedComponent_1_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( gOffloadedComponent_1_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .pcOutN_valid(  ),
       .pcOutN_bits_request(  ),
       .pcOutN_bits_moduleId(  ),
       .pcOutN_bits_portId(  ),
       .pcOutN_bits_pcValue(  ),
       .pcOutN_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_1_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_1_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_1_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_1_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_1_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_1_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_1_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_1_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_1_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_1_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_1_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_1_tag ));
  RRDistributorComponent inputDist(.clk(clk), .reset(reset),
       .io_out_0_ready( gOffloadedComponent_io_in_ready ),
       .io_out_0_valid( inputDist_io_out_0_valid ),
       .io_out_0_bits_done( inputDist_io_out_0_bits_done ),
       .io_out_0_bits_startPageId( inputDist_io_out_0_bits_startPageId ),
       .io_out_0_bits_length( inputDist_io_out_0_bits_length ),
       .io_out_0_tag( inputDist_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_in_ready ),
       .io_out_1_valid( inputDist_io_out_1_valid ),
       .io_out_1_bits_done( inputDist_io_out_1_bits_done ),
       .io_out_1_bits_startPageId( inputDist_io_out_1_bits_startPageId ),
       .io_out_1_bits_length( inputDist_io_out_1_bits_length ),
       .io_out_1_tag( inputDist_io_out_1_tag ),
       .io_in_ready( inputDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
  RRAggregatorComponent outputArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( outputArb_io_out_valid ),
       .io_out_bits_done( outputArb_io_out_bits_done ),
       .io_out_bits_pageId( outputArb_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( outputArb_io_out_tag ),
       .io_in_0_ready( outputArb_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_out_valid ),
       .io_in_0_bits_done( gOffloadedComponent_io_out_bits_done ),
       .io_in_0_bits_pageId( gOffloadedComponent_io_out_bits_pageId ),
       .io_in_0_bits_rankUpdate(  ),
       .io_in_0_tag( gOffloadedComponent_io_out_tag ),
       .io_in_1_ready( outputArb_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_out_valid ),
       .io_in_1_bits_done( gOffloadedComponent_1_io_out_bits_done ),
       .io_in_1_bits_pageId( gOffloadedComponent_1_io_out_bits_pageId ),
       .io_in_1_bits_rankUpdate(  ),
       .io_in_1_tag( gOffloadedComponent_1_io_out_tag ),
       .io_chosen(  ));
  gTaggedRRArbiter gTaggedRRArbiter(.clk(clk), .reset(reset),
       .io_out_ready( mainOff_mem_req_ready ),
       .io_out_valid( gTaggedRRArbiter_io_out_valid ),
       .io_out_bits_addr( gTaggedRRArbiter_io_out_bits_addr ),
       .io_out_bits_rw( gTaggedRRArbiter_io_out_bits_rw ),
       .io_out_bits_cached( gTaggedRRArbiter_io_out_bits_cached ),
       .io_out_bits_data( gTaggedRRArbiter_io_out_bits_data ),
       .io_out_bits_size( gTaggedRRArbiter_io_out_bits_size ),
       .io_out_tag( gTaggedRRArbiter_io_out_tag ),
       .io_in_0_ready( gTaggedRRArbiter_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_off_mem_req_valid ),
       .io_in_0_bits_addr( gOffloadedComponent_io_off_mem_req_bits_addr ),
       .io_in_0_bits_rw( gOffloadedComponent_io_off_mem_req_bits_rw ),
       .io_in_0_bits_cached( gOffloadedComponent_io_off_mem_req_bits_cached ),
       .io_in_0_bits_data( gOffloadedComponent_io_off_mem_req_bits_data ),
       .io_in_0_bits_size( gOffloadedComponent_io_off_mem_req_bits_size ),
       .io_in_0_tag( gOffloadedComponent_io_off_mem_req_tag ),
       .io_in_1_ready( gTaggedRRArbiter_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_off_mem_req_valid ),
       .io_in_1_bits_addr( gOffloadedComponent_1_io_off_mem_req_bits_addr ),
       .io_in_1_bits_rw( gOffloadedComponent_1_io_off_mem_req_bits_rw ),
       .io_in_1_bits_cached( gOffloadedComponent_1_io_off_mem_req_bits_cached ),
       .io_in_1_bits_data( gOffloadedComponent_1_io_off_mem_req_bits_data ),
       .io_in_1_bits_size( gOffloadedComponent_1_io_off_mem_req_bits_size ),
       .io_in_1_tag( gOffloadedComponent_1_io_off_mem_req_tag ),
       .io_chosen(  ));
  gTaggedDistributor gTaggedDistributor(
       .io_out_0_ready( gOffloadedComponent_io_off_mem_rep_ready ),
       .io_out_0_valid( gTaggedDistributor_io_out_0_valid ),
       .io_out_0_bits_data( gTaggedDistributor_io_out_0_bits_data ),
       .io_out_0_tag( gTaggedDistributor_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_off_mem_rep_ready ),
       .io_out_1_valid( gTaggedDistributor_io_out_1_valid ),
       .io_out_1_bits_data( gTaggedDistributor_io_out_1_bits_data ),
       .io_out_1_tag( gTaggedDistributor_io_out_1_tag ),
       .io_in_ready( gTaggedDistributor_io_in_ready ),
       .io_in_valid( mainOff_mem_rep_valid ),
       .io_in_bits_data( mainOff_mem_rep_bits_data ),
       .io_in_tag( mainOff_mem_rep_tag ),
       .io_chosen(  ));
endmodule

module RREncode_14(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_15(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_16(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module cache(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_cacheMissPipe_req_ready,
    output mainOff_cacheMissPipe_req_valid,
    output[31:0] mainOff_cacheMissPipe_req_bits,
    output[9:0] mainOff_cacheMissPipe_req_tag,
    output mainOff_cacheMissPipe_rep_ready,
    input  mainOff_cacheMissPipe_rep_valid,
    input [31:0] mainOff_cacheMissPipe_rep_bits,
    input [9:0] mainOff_cacheMissPipe_rep_tag,
    input  mainOff_dram_req_ready,
    output mainOff_dram_req_valid,
    output[31:0] mainOff_dram_req_bits_addr,
    output mainOff_dram_req_bits_rw,
    output mainOff_dram_req_bits_cached,
    output[127:0] mainOff_dram_req_bits_data,
    output[3:0] mainOff_dram_req_bits_size,
    output[9:0] mainOff_dram_req_tag,
    output mainOff_dram_rep_ready,
    input  mainOff_dram_rep_valid,
    input [127:0] mainOff_dram_rep_bits_data,
    input [9:0] mainOff_dram_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T6;
  reg[0:0] subStateTh_2;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T10;
  wire AllOffloadsValid_2;
  wire T11;
  wire T12;
  wire T13;
  reg[0:0] dramPortHadValidRequest_2;
  wire T14;
  wire T15;
  wire T16;
  wire dramPort_req_valid;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  reg[7:0] State_2;
  wire T24;
  wire T25;
  wire T26;
  wire[2:0] T27;
  wire[5:0] T28;
  wire T29;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire T38;
  reg[7:0] State_1;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[7:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[31:0] T59;
  wire T60;
  wire T61;
  reg[0:0] inputReg_2_rw;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire[5:0] T65;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  reg[0:0] subStateTh_1;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire AllOffloadsReady;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] dramPortHadReadyRequest;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  reg[0:0] dram_ready_received;
  wire T92;
  wire T93;
  wire dramPort_req_ready;
  wire[31:0] dramPort_req_bits_addr;
  wire[31:0] T94;
  wire[165:0] T95;
  wire[165:0] T96;
  wire[165:0] T97;
  wire[3:0] T98;
  wire[3:0] T99;
  wire[3:0] T100;
  reg[3:0] inputReg_2_size;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[127:0] T105;
  wire[127:0] T106;
  wire[127:0] T107;
  reg[127:0] outputReg_2_data;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[55:0] T113;
  wire[31:0] T114;
  wire[31:0] T115;
  wire[31:0] T116;
  reg[31:0] inputReg_2_addr;
  wire[31:0] T117;
  wire[31:0] T118;
  wire[31:0] T119;
  wire[31:0] T120;
  reg[31:0] inputReg_1_addr;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[31:0] T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire T128;
  reg[31:0] inputReg_0_addr;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire T133;
  wire[7:0] T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire[31:0] T141;
  wire[31:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[127:0] T146;
  wire[127:0] T147;
  wire[127:0] T148;
  wire[127:0] T149;
  wire[127:0] T150;
  wire[60:0] T151;
  wire[55:0] T152;
  wire[55:0] T153;
  wire[31:0] T154;
  wire[31:0] T155;
  wire[31:0] T156;
  reg[31:0] random_2;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[31:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  reg[31:0] burst_2;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire[31:0] T172;
  wire[31:0] T173;
  wire T174;
  wire[31:0] T175;
  wire[31:0] T176;
  wire[31:0] T177;
  wire[31:0] T178;
  reg[31:0] burst_1;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[31:0] T183;
  wire[31:0] T184;
  wire T185;
  wire[31:0] T186;
  wire[31:0] T187;
  reg[31:0] burst_0;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire[31:0] T192;
  wire[31:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[31:0] T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[31:0] T204;
  wire[31:0] T205;
  wire T206;
  wire[31:0] T207;
  wire[31:0] T208;
  wire[31:0] T209;
  wire[31:0] T210;
  reg[31:0] random_1;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire T217;
  wire[31:0] T218;
  wire[31:0] T219;
  reg[31:0] random_0;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[31:0] T224;
  wire[31:0] T225;
  wire T226;
  wire[127:0] T227;
  wire[31:0] T228;
  wire[127:0] T229;
  wire[127:0] T230;
  wire[127:0] T231;
  wire T232;
  reg[127:0] outputReg_1_data;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire[127:0] T238;
  wire[127:0] T239;
  wire[127:0] T240;
  wire[127:0] T241;
  wire[127:0] T242;
  wire[127:0] T243;
  wire[127:0] T244;
  wire[127:0] T245;
  wire T246;
  reg[127:0] outputReg_0_data;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire[127:0] T252;
  wire[127:0] T253;
  wire[127:0] T254;
  wire[127:0] T255;
  wire[127:0] T256;
  wire[127:0] T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  reg[3:0] inputReg_1_size;
  wire[3:0] T262;
  wire[3:0] T263;
  wire[3:0] T264;
  reg[3:0] inputReg_0_size;
  wire[3:0] T265;
  wire[127:0] T266;
  wire[127:0] T267;
  wire[127:0] T268;
  reg[127:0] inputReg_2_data;
  wire[127:0] T269;
  wire[127:0] T270;
  wire[127:0] T271;
  wire[127:0] T272;
  reg[127:0] inputReg_1_data;
  wire[127:0] T273;
  wire[127:0] T274;
  wire[127:0] T275;
  reg[127:0] inputReg_0_data;
  wire[127:0] T276;
  wire T277;
  wire T278;
  reg[0:0] inputReg_2_cached;
  wire T279;
  wire T280;
  wire T281;
  reg[0:0] inputReg_1_cached;
  wire T282;
  wire T283;
  reg[0:0] inputReg_0_cached;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  reg[0:0] inputReg_1_rw;
  wire T289;
  wire T290;
  reg[0:0] inputReg_0_rw;
  wire T291;
  wire[31:0] T292;
  wire[31:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[31:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire T300;
  wire T301;
  wire[7:0] T302;
  wire T303;
  wire dramPort_rep_ready;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire cacheMissPipePort_req_valid;
  wire T308;
  wire T309;
  wire T310;
  wire[7:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  reg[0:0] cacheMissPipe_valid_received_2;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[9:0] T321;
  wire[9:0] cacheMissPipePort_rep_tag;
  wire cacheMissPipePort_rep_ready;
  wire[9:0] cacheMissPipePort_req_tag;
  wire[9:0] T322;
  wire cacheMissPipePort_rep_valid;
  wire T323;
  wire T324;
  wire[4:0] T325;
  wire T326;
  wire T327;
  reg[0:0] cacheMissPipe_valid_received_1;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[9:0] T332;
  wire T333;
  wire T334;
  wire[4:0] T335;
  wire T336;
  reg[0:0] cacheMissPipe_valid_received_0;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire[9:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  reg[0:0] cacheMissPipePortHadReadyRequest;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  reg[0:0] cacheMissPipe_ready_received;
  wire T351;
  wire T352;
  wire cacheMissPipePort_req_ready;
  wire T353;
  wire T354;
  wire T355;
  reg[7:0] State_0;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire[7:0] T373;
  wire[7:0] T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[7:0] T378;
  wire[7:0] T379;
  wire[7:0] T380;
  wire[7:0] T381;
  wire[7:0] T382;
  wire[7:0] T383;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[7:0] T386;
  wire[7:0] T387;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T388;
  wire[7:0] T389;
  wire[7:0] T390;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T391;
  wire[7:0] T392;
  wire[7:0] T393;
  wire[7:0] T394;
  wire[7:0] T395;
  wire T396;
  reg[0:0] subStateTh_0;
  wire T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire[1:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire[31:0] T414;
  wire[31:0] T415;
  wire[31:0] T416;
  reg[31:0] cachedAddr_2;
  wire T417;
  wire T418;
  wire[31:0] T419;
  wire[31:0] T420;
  wire[31:0] ct;
  wire[31:0] T421;
  wire[31:0] T422;
  wire[31:0] T423;
  reg[31:0] cachedAddr_1;
  wire T424;
  wire[31:0] T425;
  wire[31:0] T426;
  wire[31:0] T427;
  wire[31:0] T428;
  reg[31:0] cachedAddr_0;
  wire T429;
  wire[31:0] T430;
  wire[31:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[7:0] T436;
  wire[7:0] T437;
  wire[7:0] T438;
  wire[7:0] T439;
  wire[7:0] T440;
  wire[7:0] T441;
  wire[7:0] T442;
  wire[7:0] T443;
  wire[7:0] T444;
  wire[7:0] T445;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T448;
  wire[7:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  reg[0:0] dram_valid_received_2;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[9:0] T486;
  wire[9:0] dramPort_rep_tag;
  wire[9:0] dramPort_req_tag;
  wire[9:0] T487;
  wire dramPort_rep_valid;
  wire T488;
  wire T489;
  wire[4:0] T490;
  wire T491;
  wire T492;
  reg[0:0] dram_valid_received_1;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire[9:0] T497;
  wire T498;
  wire T499;
  wire[4:0] T500;
  wire T501;
  reg[0:0] dram_valid_received_0;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire[9:0] T506;
  wire T507;
  wire T508;
  wire[4:0] T509;
  wire T510;
  wire T511;
  wire[4:0] T512;
  wire T513;
  wire T514;
  wire[4:0] T515;
  wire T516;
  wire T517;
  wire T518;
  wire[9:0] T519;
  wire T520;
  wire T521;
  reg[0:0] cacheMissPipePortHadValidRequest_2;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[4:0] T526;
  wire T527;
  wire T528;
  wire[4:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire[9:0] T533;
  wire T534;
  wire T535;
  wire AllOffloadsValid_1;
  wire T536;
  wire T537;
  wire T538;
  reg[0:0] dramPortHadValidRequest_1;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire[4:0] T543;
  wire T544;
  wire T545;
  wire[4:0] T546;
  wire T547;
  wire T548;
  wire T549;
  wire[9:0] T550;
  wire T551;
  wire T552;
  reg[0:0] cacheMissPipePortHadValidRequest_1;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire[4:0] T557;
  wire T558;
  wire T559;
  wire[4:0] T560;
  wire T561;
  wire T562;
  wire T563;
  wire[9:0] T564;
  wire T565;
  wire T566;
  wire AllOffloadsValid_0;
  wire T567;
  wire T568;
  wire T569;
  reg[0:0] dramPortHadValidRequest_0;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[4:0] T574;
  wire T575;
  wire T576;
  wire[4:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire[9:0] T581;
  wire T582;
  wire T583;
  reg[0:0] cacheMissPipePortHadValidRequest_0;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[4:0] T588;
  wire T589;
  wire T590;
  wire[4:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[9:0] T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[9:0] inputTag_2;
  wire[9:0] T607;
  wire[9:0] T608;
  wire[9:0] T609;
  wire[9:0] T610;
  reg[9:0] inputTag_1;
  wire[9:0] T611;
  wire[9:0] T612;
  wire[9:0] T613;
  reg[9:0] inputTag_0;
  wire[9:0] T614;

  assign io_out_tag = T0;
  assign T0 = T608 | T1;
  assign T1 = inputTag_2 & T2;
  assign T2 = {4'ha/* 10*/{T3}};
  assign T3 = T4[2'h2/* 2*/];
  assign T4 = T5[2'h2/* 2*/:1'h0/* 0*/];
  assign T5 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T6 = subStateTh_2 == 1'h0/* 0*/;
  assign T7 = T598 ? 1'h1/* 1*/ : T8;
  assign T8 = T9 ? 1'h0/* 0*/ : subStateTh_2;
  assign T9 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T10 = T534 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T11;
  assign T11 = T520 && T12;
  assign T12 = T516 || T13;
  assign T13 = ! dramPortHadValidRequest_2;
  assign T14 = T513 && T15;
  assign T15 = dramPortHadValidRequest_2 || T16;
  assign T16 = T511 && dramPort_req_valid;
  assign dramPort_req_valid = T17;
  assign T17 = T478 && T18;
  assign T18 = T477 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = T472 | T22;
  assign T22 = State_2 & T23;
  assign T23 = {4'h8/* 8*/{T3}};
  assign T24 = T451 || T25;
  assign T25 = T29 && T26;
  assign T26 = T27[2'h2/* 2*/];
  assign T27 = T28[2'h2/* 2*/:1'h0/* 0*/];
  assign T28 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T29 = T450 && T30;
  assign T30 = T32 == T31;
  assign T31 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T32 = T35 | T33;
  assign T33 = State_2 & T34;
  assign T34 = {4'h8/* 8*/{T26}};
  assign T35 = T448 | T36;
  assign T36 = State_1 & T37;
  assign T37 = {4'h8/* 8*/{T38}};
  assign T38 = T27[1'h1/* 1*/];
  assign T39 = T41 || T40;
  assign T40 = T29 && T38;
  assign T41 = T47 || T42;
  assign T42 = T43 && T38;
  assign T43 = T46 && T44;
  assign T44 = T32 == T45;
  assign T45 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T46 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T47 = T53 || T48;
  assign T48 = T49 && T38;
  assign T49 = T52 && T50;
  assign T50 = T32 == T51;
  assign T51 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T52 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T53 = T432 || T54;
  assign T54 = T55 && T38;
  assign T55 = T132 && T56;
  assign T56 = ! T57;
  assign T57 = T413 || T58;
  assign T58 = T59 == 32'h1/* 1*/;
  assign T59 = {31'h0/* 0*/, T60};
  assign T60 = T410 | T61;
  assign T61 = inputReg_2_rw & T26;
  assign T62 = T123 && T63;
  assign T63 = T64[2'h2/* 2*/];
  assign T64 = T65[2'h2/* 2*/:1'h0/* 0*/];
  assign T65 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T66 = T68 && T67;
  assign T67 = State_2 == 8'h0/* 0*/;
  assign T68 = subStateTh_2 == 1'h0/* 0*/;
  assign T69 = T71 && T70;
  assign T70 = State_1 == 8'h0/* 0*/;
  assign T71 = subStateTh_1 == 1'h0/* 0*/;
  assign T72 = T76 ? 1'h1/* 1*/ : T73;
  assign T73 = T74 ? 1'h0/* 0*/ : subStateTh_1;
  assign T74 = T75 == vThreadEncoder_io_chosen;
  assign T75 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T76 = T78 && T77;
  assign T77 = State_1 != 8'hff/* 255*/;
  assign T78 = T80 && T79;
  assign T79 = State_1 != 8'h0/* 0*/;
  assign T80 = AllOffloadsReady && T81;
  assign T81 = T82 == rThreadEncoder_io_chosen;
  assign T82 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign AllOffloadsReady = T83;
  assign T83 = T305 && T84;
  assign T84 = T91 || T85;
  assign T85 = T87 && T86;
  assign T86 = ! dramPort_req_valid;
  assign T87 = ! dramPortHadReadyRequest;
  assign T88 = T90 && T89;
  assign T89 = dramPortHadReadyRequest || dramPort_req_valid;
  assign T90 = ! AllOffloadsReady;
  assign T91 = dramPort_req_ready || dram_ready_received;
  assign T92 = T304 && T93;
  assign T93 = dram_ready_received || dramPort_req_ready;
  assign dramPort_req_ready = mainOff_dram_req_ready;
  assign mainOff_dram_req_valid = dramPort_req_valid;
  assign mainOff_dram_req_bits_addr = dramPort_req_bits_addr;
  assign dramPort_req_bits_addr = T94;
  assign T94 = T95[8'ha5/* 165*/:8'h86/* 134*/];
  assign T95 = T300 ? T97 : T96;
  assign T96 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T97 = {T292, T285, T277, T266, T98};
  assign T98 = T259 | T99;
  assign T99 = inputReg_2_size & T100;
  assign T100 = {3'h4/* 4*/{T3}};
  assign T101 = T62 ? io_in_bits_size : inputReg_2_size;
  assign io_out_valid = T102;
  assign T102 = T104 && T103;
  assign T103 = T21 == 8'hff/* 255*/;
  assign T104 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_data = T105;
  assign T105 = T229 | T106;
  assign T106 = outputReg_2_data & T107;
  assign T107 = {8'h80/* 128*/{T3}};
  assign T108 = T136 || T109;
  assign T109 = T110 && T26;
  assign T110 = T132 && T111;
  assign T111 = ! T112;
  assign T112 = T113 <= 56'h1000000/* 16777216*/;
  assign T113 = {24'h0/* 0*/, T114};
  assign T114 = T118 | T115;
  assign T115 = inputReg_2_addr & T116;
  assign T116 = {6'h20/* 32*/{T26}};
  assign T117 = T62 ? io_in_bits_addr : inputReg_2_addr;
  assign T118 = T126 | T119;
  assign T119 = inputReg_1_addr & T120;
  assign T120 = {6'h20/* 32*/{T38}};
  assign T121 = T123 && T122;
  assign T122 = T64[1'h1/* 1*/];
  assign T123 = T124 && io_in_valid;
  assign T124 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T121 ? io_in_bits_addr : inputReg_1_addr;
  assign T126 = inputReg_0_addr & T127;
  assign T127 = {6'h20/* 32*/{T128}};
  assign T128 = T27[1'h0/* 0*/];
  assign T129 = T123 && T130;
  assign T130 = T64[1'h0/* 0*/];
  assign T131 = T129 ? io_in_bits_addr : inputReg_0_addr;
  assign T132 = T135 && T133;
  assign T133 = T32 == T134;
  assign T134 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T135 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T136 = T144 || T137;
  assign T137 = T138 && T26;
  assign T138 = T143 && T139;
  assign T139 = ! T140;
  assign T140 = T141 == 32'h0/* 0*/;
  assign T141 = T142 & 32'h1/* 1*/;
  assign T142 = T114 >> 32'h2/* 2*/;
  assign T143 = T132 && T112;
  assign T144 = T145 && T26;
  assign T145 = T143 && T140;
  assign T146 = T109 ? T227 : T147;
  assign T147 = T137 ? T150 : T148;
  assign T148 = T144 ? T149 : outputReg_2_data;
  assign T149 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T150 = {67'h0/* 0*/, T151};
  assign T151 = T152 << 32'h5/* 5*/;
  assign T152 = 56'h1000000/* 16777216*/ + T153;
  assign T153 = {24'h0/* 0*/, T154};
  assign T154 = T208 | T155;
  assign T155 = random_2 & T156;
  assign T156 = {6'h20/* 32*/{T26}};
  assign T157 = T199 || T158;
  assign T158 = T159 && T26;
  assign T159 = T195 && T160;
  assign T160 = T161 == 32'h1/* 1*/;
  assign T161 = T176 | T162;
  assign T162 = burst_2 & T163;
  assign T163 = {6'h20/* 32*/{T26}};
  assign T164 = T169 || T165;
  assign T165 = T166 && T26;
  assign T166 = T145 && T167;
  assign T167 = ! T168;
  assign T168 = T161 == 32'h1/* 1*/;
  assign T169 = T62 || T170;
  assign T170 = T171 && T26;
  assign T171 = T145 && T168;
  assign T172 = T165 ? T175 : T173;
  assign T173 = T174 ? 32'h1/* 1*/ : burst_2;
  assign T174 = T62 || T170;
  assign T175 = T161 + 32'h1/* 1*/;
  assign T176 = T186 | T177;
  assign T177 = burst_1 & T178;
  assign T178 = {6'h20/* 32*/{T38}};
  assign T179 = T181 || T180;
  assign T180 = T166 && T38;
  assign T181 = T121 || T182;
  assign T182 = T171 && T38;
  assign T183 = T180 ? T175 : T184;
  assign T184 = T185 ? 32'h1/* 1*/ : burst_1;
  assign T185 = T121 || T182;
  assign T186 = burst_0 & T187;
  assign T187 = {6'h20/* 32*/{T128}};
  assign T188 = T190 || T189;
  assign T189 = T166 && T128;
  assign T190 = T129 || T191;
  assign T191 = T171 && T128;
  assign T192 = T189 ? T175 : T193;
  assign T193 = T194 ? 32'h1/* 1*/ : burst_0;
  assign T194 = T129 || T191;
  assign T195 = T145 && T196;
  assign T196 = ! T197;
  assign T197 = T154 == T198;
  assign T198 = {1'h0/* 0*/, 31'h2/* 2*/};
  assign T199 = T62 || T200;
  assign T200 = T201 && T26;
  assign T201 = T203 && T202;
  assign T202 = T161 == 32'h1/* 1*/;
  assign T203 = T145 && T197;
  assign T204 = T158 ? T207 : T205;
  assign T205 = T206 ? 32'h1/* 1*/ : random_2;
  assign T206 = T62 || T200;
  assign T207 = T154 + 32'h1/* 1*/;
  assign T208 = T218 | T209;
  assign T209 = random_1 & T210;
  assign T210 = {6'h20/* 32*/{T38}};
  assign T211 = T213 || T212;
  assign T212 = T159 && T38;
  assign T213 = T121 || T214;
  assign T214 = T201 && T38;
  assign T215 = T212 ? T207 : T216;
  assign T216 = T217 ? 32'h1/* 1*/ : random_1;
  assign T217 = T121 || T214;
  assign T218 = random_0 & T219;
  assign T219 = {6'h20/* 32*/{T128}};
  assign T220 = T222 || T221;
  assign T221 = T159 && T128;
  assign T222 = T129 || T223;
  assign T223 = T201 && T128;
  assign T224 = T221 ? T207 : T225;
  assign T225 = T226 ? 32'h1/* 1*/ : random_0;
  assign T226 = T129 || T223;
  assign T227 = {96'h0/* 0*/, T228};
  assign T228 = T114 + 32'h3e8/* 1000*/;
  assign T229 = T244 | T230;
  assign T230 = outputReg_1_data & T231;
  assign T231 = {8'h80/* 128*/{T232}};
  assign T232 = T4[1'h1/* 1*/];
  assign T233 = T235 || T234;
  assign T234 = T110 && T38;
  assign T235 = T237 || T236;
  assign T236 = T138 && T38;
  assign T237 = T145 && T38;
  assign T238 = T234 ? T243 : T239;
  assign T239 = T236 ? T242 : T240;
  assign T240 = T237 ? T241 : outputReg_1_data;
  assign T241 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T242 = {67'h0/* 0*/, T151};
  assign T243 = {96'h0/* 0*/, T228};
  assign T244 = outputReg_0_data & T245;
  assign T245 = {8'h80/* 128*/{T246}};
  assign T246 = T4[1'h0/* 0*/];
  assign T247 = T249 || T248;
  assign T248 = T110 && T128;
  assign T249 = T251 || T250;
  assign T250 = T138 && T128;
  assign T251 = T145 && T128;
  assign T252 = T248 ? T257 : T253;
  assign T253 = T250 ? T256 : T254;
  assign T254 = T251 ? T255 : outputReg_0_data;
  assign T255 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T256 = {67'h0/* 0*/, T151};
  assign T257 = {96'h0/* 0*/, T228};
  assign io_in_ready = T258;
  assign T258 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T259 = T263 | T260;
  assign T260 = inputReg_1_size & T261;
  assign T261 = {3'h4/* 4*/{T232}};
  assign T262 = T121 ? io_in_bits_size : inputReg_1_size;
  assign T263 = inputReg_0_size & T264;
  assign T264 = {3'h4/* 4*/{T246}};
  assign T265 = T129 ? io_in_bits_size : inputReg_0_size;
  assign T266 = T270 | T267;
  assign T267 = inputReg_2_data & T268;
  assign T268 = {8'h80/* 128*/{T3}};
  assign T269 = T62 ? io_in_bits_data : inputReg_2_data;
  assign T270 = T274 | T271;
  assign T271 = inputReg_1_data & T272;
  assign T272 = {8'h80/* 128*/{T232}};
  assign T273 = T121 ? io_in_bits_data : inputReg_1_data;
  assign T274 = inputReg_0_data & T275;
  assign T275 = {8'h80/* 128*/{T246}};
  assign T276 = T129 ? io_in_bits_data : inputReg_0_data;
  assign T277 = T280 | T278;
  assign T278 = inputReg_2_cached & T3;
  assign T279 = T62 ? io_in_bits_cached : inputReg_2_cached;
  assign T280 = T283 | T281;
  assign T281 = inputReg_1_cached & T232;
  assign T282 = T121 ? io_in_bits_cached : inputReg_1_cached;
  assign T283 = inputReg_0_cached & T246;
  assign T284 = T129 ? io_in_bits_cached : inputReg_0_cached;
  assign T285 = T287 | T286;
  assign T286 = inputReg_2_rw & T3;
  assign T287 = T290 | T288;
  assign T288 = inputReg_1_rw & T232;
  assign T289 = T121 ? io_in_bits_rw : inputReg_1_rw;
  assign T290 = inputReg_0_rw & T246;
  assign T291 = T129 ? io_in_bits_rw : inputReg_0_rw;
  assign T292 = T295 | T293;
  assign T293 = inputReg_2_addr & T294;
  assign T294 = {6'h20/* 32*/{T3}};
  assign T295 = T298 | T296;
  assign T296 = inputReg_1_addr & T297;
  assign T297 = {6'h20/* 32*/{T232}};
  assign T298 = inputReg_0_addr & T299;
  assign T299 = {6'h20/* 32*/{T246}};
  assign T300 = T303 && T301;
  assign T301 = T21 == T302;
  assign T302 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T303 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign mainOff_dram_rep_ready = dramPort_rep_ready;
  assign dramPort_rep_ready = 1'h1/* 1*/;
  assign T304 = ! AllOffloadsReady;
  assign T305 = T350 || T306;
  assign T306 = T346 && T307;
  assign T307 = ! cacheMissPipePort_req_valid;
  assign cacheMissPipePort_req_valid = T308;
  assign T308 = T313 && T309;
  assign T309 = T312 && T310;
  assign T310 = T21 == T311;
  assign T311 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T312 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T313 = T345 && T314;
  assign T314 = ! T315;
  assign T315 = T326 | T316;
  assign T316 = cacheMissPipe_valid_received_2 & T3;
  assign T317 = T323 && T318;
  assign T318 = cacheMissPipe_valid_received_2 || T319;
  assign T319 = cacheMissPipePort_rep_valid && T320;
  assign T320 = cacheMissPipePort_rep_tag == T321;
  assign T321 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign cacheMissPipePort_rep_tag = mainOff_cacheMissPipe_rep_tag;
  assign mainOff_cacheMissPipe_rep_ready = cacheMissPipePort_rep_ready;
  assign cacheMissPipePort_rep_ready = 1'h1/* 1*/;
  assign mainOff_cacheMissPipe_req_tag = cacheMissPipePort_req_tag;
  assign cacheMissPipePort_req_tag = T322;
  assign T322 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign cacheMissPipePort_rep_valid = mainOff_cacheMissPipe_rep_valid;
  assign mainOff_cacheMissPipe_req_valid = cacheMissPipePort_req_valid;
  assign T323 = ! T324;
  assign T324 = T325 == 5'h2/* 2*/;
  assign T325 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T326 = T336 | T327;
  assign T327 = cacheMissPipe_valid_received_1 & T232;
  assign T328 = T333 && T329;
  assign T329 = cacheMissPipe_valid_received_1 || T330;
  assign T330 = cacheMissPipePort_rep_valid && T331;
  assign T331 = cacheMissPipePort_rep_tag == T332;
  assign T332 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T333 = ! T334;
  assign T334 = T335 == 5'h1/* 1*/;
  assign T335 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T336 = cacheMissPipe_valid_received_0 & T246;
  assign T337 = T342 && T338;
  assign T338 = cacheMissPipe_valid_received_0 || T339;
  assign T339 = cacheMissPipePort_rep_valid && T340;
  assign T340 = cacheMissPipePort_rep_tag == T341;
  assign T341 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T346 = ! cacheMissPipePortHadReadyRequest;
  assign T347 = T349 && T348;
  assign T348 = cacheMissPipePortHadReadyRequest || cacheMissPipePort_req_valid;
  assign T349 = ! AllOffloadsReady;
  assign T350 = cacheMissPipePort_req_ready || cacheMissPipe_ready_received;
  assign T351 = T353 && T352;
  assign T352 = cacheMissPipe_ready_received || cacheMissPipePort_req_ready;
  assign cacheMissPipePort_req_ready = mainOff_cacheMissPipe_req_ready;
  assign T353 = ! AllOffloadsReady;
  assign T354 = T396 && T355;
  assign T355 = State_0 == 8'h0/* 0*/;
  assign T356 = T358 || T357;
  assign T357 = T29 && T128;
  assign T358 = T360 || T359;
  assign T359 = T43 && T128;
  assign T360 = T362 || T361;
  assign T361 = T49 && T128;
  assign T362 = T364 || T363;
  assign T363 = T55 && T128;
  assign T364 = T367 || T365;
  assign T365 = T366 && T128;
  assign T366 = T132 && T57;
  assign T367 = T129 || T368;
  assign T368 = T369 && T246;
  assign T369 = T370 && io_out_ready;
  assign T370 = T372 && T371;
  assign T371 = T21 == 8'hff/* 255*/;
  assign T372 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T373 = T357 ? 8'hff/* 255*/ : T374;
  assign T374 = T359 ? T395 : T375;
  assign T375 = T361 ? T394 : T376;
  assign T376 = T363 ? T393 : T377;
  assign T377 = T365 ? T392 : T378;
  assign T378 = T368 ? T381 : T379;
  assign T379 = T129 ? T380 : State_0;
  assign T380 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T381 = T385 | T382;
  assign T382 = EmitReturnState_2 & T383;
  assign T383 = {4'h8/* 8*/{T3}};
  assign T384 = T25 ? 8'h0/* 0*/ : EmitReturnState_2;
  assign T385 = T389 | T386;
  assign T386 = EmitReturnState_1 & T387;
  assign T387 = {4'h8/* 8*/{T232}};
  assign T388 = T40 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T389 = EmitReturnState_0 & T390;
  assign T390 = {4'h8/* 8*/{T246}};
  assign T391 = T357 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T392 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T393 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T394 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T395 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T396 = subStateTh_0 == 1'h0/* 0*/;
  assign T397 = T401 ? 1'h1/* 1*/ : T398;
  assign T398 = T399 ? 1'h0/* 0*/ : subStateTh_0;
  assign T399 = T400 == vThreadEncoder_io_chosen;
  assign T400 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T401 = T403 && T402;
  assign T402 = State_0 != 8'hff/* 255*/;
  assign T403 = T405 && T404;
  assign T404 = State_0 != 8'h0/* 0*/;
  assign T405 = AllOffloadsReady && T406;
  assign T406 = T407 == rThreadEncoder_io_chosen;
  assign T407 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T408 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T409 = T62 ? io_in_bits_rw : inputReg_2_rw;
  assign T410 = T412 | T411;
  assign T411 = inputReg_1_rw & T38;
  assign T412 = inputReg_0_rw & T128;
  assign T413 = ct == T414;
  assign T414 = T421 | T415;
  assign T415 = cachedAddr_2 & T416;
  assign T416 = {6'h20/* 32*/{T26}};
  assign T417 = T62 || T418;
  assign T418 = T55 && T26;
  assign T419 = T418 ? ct : T420;
  assign T420 = T62 ? 32'h0/* 0*/ : cachedAddr_2;
  assign ct = T114 >> 32'h4/* 4*/;
  assign T421 = T427 | T422;
  assign T422 = cachedAddr_1 & T423;
  assign T423 = {6'h20/* 32*/{T38}};
  assign T424 = T121 || T54;
  assign T425 = T54 ? ct : T426;
  assign T426 = T121 ? 32'h0/* 0*/ : cachedAddr_1;
  assign T427 = cachedAddr_0 & T428;
  assign T428 = {6'h20/* 32*/{T128}};
  assign T429 = T129 || T363;
  assign T430 = T363 ? ct : T431;
  assign T431 = T129 ? 32'h0/* 0*/ : cachedAddr_0;
  assign T432 = T434 || T433;
  assign T433 = T366 && T38;
  assign T434 = T121 || T435;
  assign T435 = T369 && T232;
  assign T436 = T40 ? 8'hff/* 255*/ : T437;
  assign T437 = T42 ? T447 : T438;
  assign T438 = T48 ? T446 : T439;
  assign T439 = T54 ? T445 : T440;
  assign T440 = T433 ? T444 : T441;
  assign T441 = T435 ? T381 : T442;
  assign T442 = T121 ? T443 : State_1;
  assign T443 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T444 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T445 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T446 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T447 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T448 = State_0 & T449;
  assign T449 = {4'h8/* 8*/{T128}};
  assign T450 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T451 = T453 || T452;
  assign T452 = T43 && T26;
  assign T453 = T455 || T454;
  assign T454 = T49 && T26;
  assign T455 = T456 || T418;
  assign T456 = T458 || T457;
  assign T457 = T366 && T26;
  assign T458 = T62 || T459;
  assign T459 = T369 && T3;
  assign T460 = T25 ? 8'hff/* 255*/ : T461;
  assign T461 = T452 ? T471 : T462;
  assign T462 = T454 ? T470 : T463;
  assign T463 = T418 ? T469 : T464;
  assign T464 = T457 ? T468 : T465;
  assign T465 = T459 ? T381 : T466;
  assign T466 = T62 ? T467 : State_2;
  assign T467 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T468 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T469 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T470 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T471 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T472 = T475 | T473;
  assign T473 = State_1 & T474;
  assign T474 = {4'h8/* 8*/{T232}};
  assign T475 = State_0 & T476;
  assign T476 = {4'h8/* 8*/{T246}};
  assign T477 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T478 = T510 && T479;
  assign T479 = ! T480;
  assign T480 = T491 | T481;
  assign T481 = dram_valid_received_2 & T3;
  assign T482 = T488 && T483;
  assign T483 = dram_valid_received_2 || T484;
  assign T484 = dramPort_rep_valid && T485;
  assign T485 = dramPort_rep_tag == T486;
  assign T486 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign dramPort_rep_tag = mainOff_dram_rep_tag;
  assign mainOff_dram_req_tag = dramPort_req_tag;
  assign dramPort_req_tag = T487;
  assign T487 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramPort_rep_valid = mainOff_dram_rep_valid;
  assign T488 = ! T489;
  assign T489 = T490 == 5'h2/* 2*/;
  assign T490 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T491 = T501 | T492;
  assign T492 = dram_valid_received_1 & T232;
  assign T493 = T498 && T494;
  assign T494 = dram_valid_received_1 || T495;
  assign T495 = dramPort_rep_valid && T496;
  assign T496 = dramPort_rep_tag == T497;
  assign T497 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T498 = ! T499;
  assign T499 = T500 == 5'h1/* 1*/;
  assign T500 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T501 = dram_valid_received_0 & T246;
  assign T502 = T507 && T503;
  assign T503 = dram_valid_received_0 || T504;
  assign T504 = dramPort_rep_valid && T505;
  assign T505 = dramPort_rep_tag == T506;
  assign T506 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T507 = ! T508;
  assign T508 = T509 == 5'h0/* 0*/;
  assign T509 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T510 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T511 = 5'h2/* 2*/ == T512;
  assign T512 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T513 = ! T514;
  assign T514 = T515 == 5'h2/* 2*/;
  assign T515 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T516 = T517 || dram_valid_received_2;
  assign T517 = dramPort_rep_valid && T518;
  assign T518 = dramPort_rep_tag == T519;
  assign T519 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T520 = T530 || T521;
  assign T521 = ! cacheMissPipePortHadValidRequest_2;
  assign T522 = T527 && T523;
  assign T523 = cacheMissPipePortHadValidRequest_2 || T524;
  assign T524 = T525 && cacheMissPipePort_req_valid;
  assign T525 = 5'h2/* 2*/ == T526;
  assign T526 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T527 = ! T528;
  assign T528 = T529 == 5'h2/* 2*/;
  assign T529 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T530 = T531 || cacheMissPipe_valid_received_2;
  assign T531 = cacheMissPipePort_rep_valid && T532;
  assign T532 = cacheMissPipePort_rep_tag == T533;
  assign T533 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T534 = subStateTh_2 == 1'h1/* 1*/;
  assign T535 = T565 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T536;
  assign T536 = T551 && T537;
  assign T537 = T547 || T538;
  assign T538 = ! dramPortHadValidRequest_1;
  assign T539 = T544 && T540;
  assign T540 = dramPortHadValidRequest_1 || T541;
  assign T541 = T542 && dramPort_req_valid;
  assign T542 = 5'h1/* 1*/ == T543;
  assign T543 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T544 = ! T545;
  assign T545 = T546 == 5'h1/* 1*/;
  assign T546 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T547 = T548 || dram_valid_received_1;
  assign T548 = dramPort_rep_valid && T549;
  assign T549 = dramPort_rep_tag == T550;
  assign T550 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T551 = T561 || T552;
  assign T552 = ! cacheMissPipePortHadValidRequest_1;
  assign T553 = T558 && T554;
  assign T554 = cacheMissPipePortHadValidRequest_1 || T555;
  assign T555 = T556 && cacheMissPipePort_req_valid;
  assign T556 = 5'h1/* 1*/ == T557;
  assign T557 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T558 = ! T559;
  assign T559 = T560 == 5'h1/* 1*/;
  assign T560 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T561 = T562 || cacheMissPipe_valid_received_1;
  assign T562 = cacheMissPipePort_rep_valid && T563;
  assign T563 = cacheMissPipePort_rep_tag == T564;
  assign T564 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T565 = subStateTh_1 == 1'h1/* 1*/;
  assign T566 = T596 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T567;
  assign T567 = T582 && T568;
  assign T568 = T578 || T569;
  assign T569 = ! dramPortHadValidRequest_0;
  assign T570 = T575 && T571;
  assign T571 = dramPortHadValidRequest_0 || T572;
  assign T572 = T573 && dramPort_req_valid;
  assign T573 = 5'h0/* 0*/ == T574;
  assign T574 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T575 = ! T576;
  assign T576 = T577 == 5'h0/* 0*/;
  assign T577 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T578 = T579 || dram_valid_received_0;
  assign T579 = dramPort_rep_valid && T580;
  assign T580 = dramPort_rep_tag == T581;
  assign T581 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T582 = T592 || T583;
  assign T583 = ! cacheMissPipePortHadValidRequest_0;
  assign T584 = T589 && T585;
  assign T585 = cacheMissPipePortHadValidRequest_0 || T586;
  assign T586 = T587 && cacheMissPipePort_req_valid;
  assign T587 = 5'h0/* 0*/ == T588;
  assign T588 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T589 = ! T590;
  assign T590 = T591 == 5'h0/* 0*/;
  assign T591 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T592 = T593 || cacheMissPipe_valid_received_0;
  assign T593 = cacheMissPipePort_rep_valid && T594;
  assign T594 = cacheMissPipePort_rep_tag == T595;
  assign T595 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T596 = subStateTh_0 == 1'h1/* 1*/;
  assign T597 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T598 = T600 && T599;
  assign T599 = State_2 != 8'hff/* 255*/;
  assign T600 = T602 && T601;
  assign T601 = State_2 != 8'h0/* 0*/;
  assign T602 = AllOffloadsReady && T603;
  assign T603 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign T604 = subStateTh_1 == 1'h0/* 0*/;
  assign T605 = subStateTh_0 == 1'h0/* 0*/;
  assign T606 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T607 = T62 ? io_in_tag : inputTag_2;
  assign T608 = T612 | T609;
  assign T609 = inputTag_1 & T610;
  assign T610 = {4'ha/* 10*/{T232}};
  assign T611 = T121 ? io_in_tag : inputTag_1;
  assign T612 = inputTag_0 & T613;
  assign T613 = {4'ha/* 10*/{T246}};
  assign T614 = T129 ? io_in_tag : inputTag_0;
  RREncode_14 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T605 ),
       .io_valid_1( T604 ),
       .io_valid_2( T6 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T606 ));
  RREncode_15 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T566 ),
       .io_valid_1( T535 ),
       .io_valid_2( T10 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T597 ));
  RREncode_16 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T354 ),
       .io_valid_1( T69 ),
       .io_valid_2( T66 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T408 ));

  always @(posedge clk) begin
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T7;
    dramPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T14;
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T24) begin
      State_2 <= T460;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T39) begin
      State_1 <= T436;
    end
    if(T62) begin
      inputReg_2_rw <= T409;
    end
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T72;
    dramPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T88;
    dram_ready_received <= reset ? 1'h0/* 0*/ : T92;
    if(T62) begin
      inputReg_2_size <= T101;
    end
    if(T108) begin
      outputReg_2_data <= T146;
    end
    if(T62) begin
      inputReg_2_addr <= T117;
    end
    if(T121) begin
      inputReg_1_addr <= T125;
    end
    if(T129) begin
      inputReg_0_addr <= T131;
    end
    if(reset) begin
      random_2 <= 32'h1/* 1*/;
    end else if(T157) begin
      random_2 <= T204;
    end
    if(reset) begin
      burst_2 <= 32'h1/* 1*/;
    end else if(T164) begin
      burst_2 <= T172;
    end
    if(reset) begin
      burst_1 <= 32'h1/* 1*/;
    end else if(T179) begin
      burst_1 <= T183;
    end
    if(reset) begin
      burst_0 <= 32'h1/* 1*/;
    end else if(T188) begin
      burst_0 <= T192;
    end
    if(reset) begin
      random_1 <= 32'h1/* 1*/;
    end else if(T211) begin
      random_1 <= T215;
    end
    if(reset) begin
      random_0 <= 32'h1/* 1*/;
    end else if(T220) begin
      random_0 <= T224;
    end
    if(T233) begin
      outputReg_1_data <= T238;
    end
    if(T247) begin
      outputReg_0_data <= T252;
    end
    if(T121) begin
      inputReg_1_size <= T262;
    end
    if(T129) begin
      inputReg_0_size <= T265;
    end
    if(T62) begin
      inputReg_2_data <= T269;
    end
    if(T121) begin
      inputReg_1_data <= T273;
    end
    if(T129) begin
      inputReg_0_data <= T276;
    end
    if(T62) begin
      inputReg_2_cached <= T279;
    end
    if(T121) begin
      inputReg_1_cached <= T282;
    end
    if(T129) begin
      inputReg_0_cached <= T284;
    end
    if(T121) begin
      inputReg_1_rw <= T289;
    end
    if(T129) begin
      inputReg_0_rw <= T291;
    end
    cacheMissPipe_valid_received_2 <= reset ? 1'h0/* 0*/ : T317;
    cacheMissPipe_valid_received_1 <= reset ? 1'h0/* 0*/ : T328;
    cacheMissPipe_valid_received_0 <= reset ? 1'h0/* 0*/ : T337;
    cacheMissPipePortHadReadyRequest <= reset ? 1'h0/* 0*/ : T347;
    cacheMissPipe_ready_received <= reset ? 1'h0/* 0*/ : T351;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T356) begin
      State_0 <= T373;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T25) begin
      EmitReturnState_2 <= T384;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T40) begin
      EmitReturnState_1 <= T388;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T357) begin
      EmitReturnState_0 <= T391;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T397;
    if(reset) begin
      cachedAddr_2 <= 32'h0/* 0*/;
    end else if(T417) begin
      cachedAddr_2 <= T419;
    end
    if(reset) begin
      cachedAddr_1 <= 32'h0/* 0*/;
    end else if(T424) begin
      cachedAddr_1 <= T425;
    end
    if(reset) begin
      cachedAddr_0 <= 32'h0/* 0*/;
    end else if(T429) begin
      cachedAddr_0 <= T430;
    end
    dram_valid_received_2 <= reset ? 1'h0/* 0*/ : T482;
    dram_valid_received_1 <= reset ? 1'h0/* 0*/ : T493;
    dram_valid_received_0 <= reset ? 1'h0/* 0*/ : T502;
    cacheMissPipePortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T522;
    dramPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T539;
    cacheMissPipePortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T553;
    dramPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T570;
    cacheMissPipePortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T584;
    if(T62) begin
      inputTag_2 <= T607;
    end
    if(T121) begin
      inputTag_1 <= T611;
    end
    if(T129) begin
      inputTag_0 <= T614;
    end
  end
endmodule

module gPipe_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_1};
  assign io_out_valid = valids_1;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module gOffloadedComponent_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dram_req_ready,
    output mainOff_dram_req_valid,
    output[31:0] mainOff_dram_req_bits_addr,
    output mainOff_dram_req_bits_rw,
    output mainOff_dram_req_bits_cached,
    output[127:0] mainOff_dram_req_bits_data,
    output[3:0] mainOff_dram_req_bits_size,
    output[9:0] mainOff_dram_req_tag,
    output mainOff_dram_rep_ready,
    input  mainOff_dram_rep_valid,
    input [127:0] mainOff_dram_rep_bits_data,
    input [9:0] mainOff_dram_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_dram_req_valid;
  wire[31:0] mainComp_mainOff_dram_req_bits_addr;
  wire mainComp_io_out_valid;
  wire[127:0] mainComp_io_out_bits_data;
  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dram_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_cacheMissPipe_rep_ready;
  wire[9:0] mainComp_mainOff_cacheMissPipe_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_cacheMissPipe_req_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dram_req_tag;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_dram_req_valid = mainComp_mainOff_dram_req_valid;
  assign mainOff_dram_req_bits_addr = mainComp_mainOff_dram_req_bits_addr;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_data = mainComp_io_out_bits_data;
  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dram_rep_ready = mainComp_mainOff_dram_rep_ready;
  assign mainOff_dram_req_tag = mainComp_mainOff_dram_req_tag;
  cache mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data( mainComp_io_out_bits_data ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_cacheMissPipe_req_ready( offComp_io_in_ready ),
       .mainOff_cacheMissPipe_req_valid( mainComp_mainOff_cacheMissPipe_req_valid ),
       .mainOff_cacheMissPipe_req_bits(  ),
       .mainOff_cacheMissPipe_req_tag( mainComp_mainOff_cacheMissPipe_req_tag ),
       .mainOff_cacheMissPipe_rep_ready( mainComp_mainOff_cacheMissPipe_rep_ready ),
       .mainOff_cacheMissPipe_rep_valid( offComp_io_out_valid ),
       .mainOff_cacheMissPipe_rep_bits(  ),
       .mainOff_cacheMissPipe_rep_tag( offComp_io_out_tag ),
       .mainOff_dram_req_ready( mainOff_dram_req_ready ),
       .mainOff_dram_req_valid( mainComp_mainOff_dram_req_valid ),
       .mainOff_dram_req_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .mainOff_dram_req_bits_rw(  ),
       .mainOff_dram_req_bits_cached(  ),
       .mainOff_dram_req_bits_data(  ),
       .mainOff_dram_req_bits_size(  ),
       .mainOff_dram_req_tag( mainComp_mainOff_dram_req_tag ),
       .mainOff_dram_rep_ready( mainComp_mainOff_dram_rep_ready ),
       .mainOff_dram_rep_valid( mainOff_dram_rep_valid ),
       .mainOff_dram_rep_bits_data(  ),
       .mainOff_dram_rep_tag( mainOff_dram_rep_tag ));
  gPipe_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_cacheMissPipe_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_cacheMissPipe_req_tag ),
       .io_out_ready( mainComp_mainOff_cacheMissPipe_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_17(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module RREncode_18(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module RREncode_19(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module dram(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank0_req_ready,
    output mainOff_dramBank0_req_valid,
    output[31:0] mainOff_dramBank0_req_bits,
    output[9:0] mainOff_dramBank0_req_tag,
    output mainOff_dramBank0_rep_ready,
    input  mainOff_dramBank0_rep_valid,
    input [31:0] mainOff_dramBank0_rep_bits,
    input [9:0] mainOff_dramBank0_rep_tag,
    input  mainOff_dramBank1_req_ready,
    output mainOff_dramBank1_req_valid,
    output[31:0] mainOff_dramBank1_req_bits,
    output[9:0] mainOff_dramBank1_req_tag,
    output mainOff_dramBank1_rep_ready,
    input  mainOff_dramBank1_rep_valid,
    input [31:0] mainOff_dramBank1_rep_bits,
    input [9:0] mainOff_dramBank1_rep_tag,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire T0;
  wire[3:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_7;
  wire T3;
  wire T4;
  wire T5;
  wire[7:0] T6;
  wire[22:0] T7;
  wire[3:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_7;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] dramBank7PortHadValidRequest_7;
  wire T12;
  wire T13;
  wire T14;
  wire dramBank7Port_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire[7:0] T23;
  wire[22:0] T24;
  wire[3:0] rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_7;
  wire T26;
  wire T27;
  wire T28;
  wire[3:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire AllOffloadsReady;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg[0:0] dramBank7PortHadReadyRequest;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg[0:0] dramBank7_ready_received;
  wire T46;
  wire T47;
  wire dramBank7Port_req_ready;
  wire dramBank7Port_rep_ready;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire dramBank6Port_req_valid;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  reg[0:0] dramBank6_valid_received_7;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[9:0] T66;
  wire[9:0] dramBank6Port_rep_tag;
  wire dramBank6Port_rep_ready;
  wire[9:0] dramBank6Port_req_tag;
  wire[9:0] T67;
  wire dramBank6Port_rep_valid;
  wire T68;
  wire T69;
  wire[4:0] T70;
  wire T71;
  wire T72;
  wire T73;
  reg[0:0] dramBank6_valid_received_6;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[9:0] T78;
  wire T79;
  wire T80;
  wire[4:0] T81;
  wire T82;
  wire T83;
  wire T84;
  reg[0:0] dramBank6_valid_received_5;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[9:0] T89;
  wire T90;
  wire T91;
  wire[4:0] T92;
  wire T93;
  wire T94;
  wire T95;
  reg[0:0] dramBank6_valid_received_4;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[9:0] T100;
  wire T101;
  wire T102;
  wire[4:0] T103;
  wire T104;
  wire T105;
  wire T106;
  reg[0:0] dramBank6_valid_received_3;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[9:0] T111;
  wire T112;
  wire T113;
  wire[4:0] T114;
  wire T115;
  wire T116;
  wire T117;
  reg[0:0] dramBank6_valid_received_2;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[9:0] T122;
  wire T123;
  wire T124;
  wire[4:0] T125;
  wire T126;
  wire T127;
  wire T128;
  reg[0:0] dramBank6_valid_received_1;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[9:0] T133;
  wire T134;
  wire T135;
  wire[4:0] T136;
  wire T137;
  wire T138;
  reg[0:0] dramBank6_valid_received_0;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[9:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  reg[0:0] dramBank6PortHadReadyRequest;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] dramBank6_ready_received;
  wire T153;
  wire T154;
  wire dramBank6Port_req_ready;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire dramBank5Port_req_valid;
  wire T160;
  wire T161;
  wire T162;
  wire[7:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  reg[0:0] dramBank5_valid_received_7;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[9:0] T173;
  wire[9:0] dramBank5Port_rep_tag;
  wire dramBank5Port_rep_ready;
  wire[9:0] dramBank5Port_req_tag;
  wire[9:0] T174;
  wire dramBank5Port_rep_valid;
  wire T175;
  wire T176;
  wire[4:0] T177;
  wire T178;
  wire T179;
  reg[0:0] dramBank5_valid_received_6;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[9:0] T184;
  wire T185;
  wire T186;
  wire[4:0] T187;
  wire T188;
  wire T189;
  reg[0:0] dramBank5_valid_received_5;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[9:0] T194;
  wire T195;
  wire T196;
  wire[4:0] T197;
  wire T198;
  wire T199;
  reg[0:0] dramBank5_valid_received_4;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[9:0] T204;
  wire T205;
  wire T206;
  wire[4:0] T207;
  wire T208;
  wire T209;
  reg[0:0] dramBank5_valid_received_3;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[9:0] T214;
  wire T215;
  wire T216;
  wire[4:0] T217;
  wire T218;
  wire T219;
  reg[0:0] dramBank5_valid_received_2;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[9:0] T224;
  wire T225;
  wire T226;
  wire[4:0] T227;
  wire T228;
  wire T229;
  reg[0:0] dramBank5_valid_received_1;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire[9:0] T234;
  wire T235;
  wire T236;
  wire[4:0] T237;
  wire T238;
  reg[0:0] dramBank5_valid_received_0;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire[9:0] T243;
  wire T244;
  wire T245;
  wire[4:0] T246;
  wire T247;
  wire T248;
  reg[0:0] dramBank5PortHadReadyRequest;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] dramBank5_ready_received;
  wire T253;
  wire T254;
  wire dramBank5Port_req_ready;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire dramBank4Port_req_valid;
  wire T260;
  wire T261;
  wire T262;
  wire[7:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  reg[0:0] dramBank4_valid_received_7;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[9:0] T273;
  wire[9:0] dramBank4Port_rep_tag;
  wire dramBank4Port_rep_ready;
  wire[9:0] dramBank4Port_req_tag;
  wire[9:0] T274;
  wire dramBank4Port_rep_valid;
  wire T275;
  wire T276;
  wire[4:0] T277;
  wire T278;
  wire T279;
  reg[0:0] dramBank4_valid_received_6;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[9:0] T284;
  wire T285;
  wire T286;
  wire[4:0] T287;
  wire T288;
  wire T289;
  reg[0:0] dramBank4_valid_received_5;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[9:0] T294;
  wire T295;
  wire T296;
  wire[4:0] T297;
  wire T298;
  wire T299;
  reg[0:0] dramBank4_valid_received_4;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[9:0] T304;
  wire T305;
  wire T306;
  wire[4:0] T307;
  wire T308;
  wire T309;
  reg[0:0] dramBank4_valid_received_3;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire[9:0] T314;
  wire T315;
  wire T316;
  wire[4:0] T317;
  wire T318;
  wire T319;
  reg[0:0] dramBank4_valid_received_2;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[9:0] T324;
  wire T325;
  wire T326;
  wire[4:0] T327;
  wire T328;
  wire T329;
  reg[0:0] dramBank4_valid_received_1;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire T335;
  wire T336;
  wire[4:0] T337;
  wire T338;
  reg[0:0] dramBank4_valid_received_0;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire[9:0] T343;
  wire T344;
  wire T345;
  wire[4:0] T346;
  wire T347;
  wire T348;
  reg[0:0] dramBank4PortHadReadyRequest;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  reg[0:0] dramBank4_ready_received;
  wire T353;
  wire T354;
  wire dramBank4Port_req_ready;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire dramBank3Port_req_valid;
  wire T360;
  wire T361;
  wire T362;
  wire[7:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  reg[0:0] dramBank3_valid_received_7;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire[9:0] T373;
  wire[9:0] dramBank3Port_rep_tag;
  wire dramBank3Port_rep_ready;
  wire[9:0] dramBank3Port_req_tag;
  wire[9:0] T374;
  wire dramBank3Port_rep_valid;
  wire T375;
  wire T376;
  wire[4:0] T377;
  wire T378;
  wire T379;
  reg[0:0] dramBank3_valid_received_6;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire[9:0] T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire T388;
  wire T389;
  reg[0:0] dramBank3_valid_received_5;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[9:0] T394;
  wire T395;
  wire T396;
  wire[4:0] T397;
  wire T398;
  wire T399;
  reg[0:0] dramBank3_valid_received_4;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[9:0] T404;
  wire T405;
  wire T406;
  wire[4:0] T407;
  wire T408;
  wire T409;
  reg[0:0] dramBank3_valid_received_3;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire[9:0] T414;
  wire T415;
  wire T416;
  wire[4:0] T417;
  wire T418;
  wire T419;
  reg[0:0] dramBank3_valid_received_2;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[9:0] T424;
  wire T425;
  wire T426;
  wire[4:0] T427;
  wire T428;
  wire T429;
  reg[0:0] dramBank3_valid_received_1;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire[9:0] T434;
  wire T435;
  wire T436;
  wire[4:0] T437;
  wire T438;
  reg[0:0] dramBank3_valid_received_0;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire[9:0] T443;
  wire T444;
  wire T445;
  wire[4:0] T446;
  wire T447;
  wire T448;
  reg[0:0] dramBank3PortHadReadyRequest;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] dramBank3_ready_received;
  wire T453;
  wire T454;
  wire dramBank3Port_req_ready;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire dramBank2Port_req_valid;
  wire T460;
  wire T461;
  wire T462;
  wire[7:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] dramBank2_valid_received_7;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire[9:0] T473;
  wire[9:0] dramBank2Port_rep_tag;
  wire dramBank2Port_rep_ready;
  wire[9:0] dramBank2Port_req_tag;
  wire[9:0] T474;
  wire dramBank2Port_rep_valid;
  wire T475;
  wire T476;
  wire[4:0] T477;
  wire T478;
  wire T479;
  reg[0:0] dramBank2_valid_received_6;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[9:0] T484;
  wire T485;
  wire T486;
  wire[4:0] T487;
  wire T488;
  wire T489;
  reg[0:0] dramBank2_valid_received_5;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[9:0] T494;
  wire T495;
  wire T496;
  wire[4:0] T497;
  wire T498;
  wire T499;
  reg[0:0] dramBank2_valid_received_4;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[9:0] T504;
  wire T505;
  wire T506;
  wire[4:0] T507;
  wire T508;
  wire T509;
  reg[0:0] dramBank2_valid_received_3;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire[9:0] T514;
  wire T515;
  wire T516;
  wire[4:0] T517;
  wire T518;
  wire T519;
  reg[0:0] dramBank2_valid_received_2;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[9:0] T524;
  wire T525;
  wire T526;
  wire[4:0] T527;
  wire T528;
  wire T529;
  reg[0:0] dramBank2_valid_received_1;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[9:0] T534;
  wire T535;
  wire T536;
  wire[4:0] T537;
  wire T538;
  reg[0:0] dramBank2_valid_received_0;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire[9:0] T543;
  wire T544;
  wire T545;
  wire[4:0] T546;
  wire T547;
  wire T548;
  reg[0:0] dramBank2PortHadReadyRequest;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  reg[0:0] dramBank2_ready_received;
  wire T553;
  wire T554;
  wire dramBank2Port_req_ready;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire dramBank1Port_req_valid;
  wire T560;
  wire T561;
  wire T562;
  wire[7:0] T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  reg[0:0] dramBank1_valid_received_7;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire[9:0] T573;
  wire[9:0] dramBank1Port_rep_tag;
  wire dramBank1Port_rep_ready;
  wire[9:0] dramBank1Port_req_tag;
  wire[9:0] T574;
  wire dramBank1Port_rep_valid;
  wire T575;
  wire T576;
  wire[4:0] T577;
  wire T578;
  wire T579;
  reg[0:0] dramBank1_valid_received_6;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire[9:0] T584;
  wire T585;
  wire T586;
  wire[4:0] T587;
  wire T588;
  wire T589;
  reg[0:0] dramBank1_valid_received_5;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire[9:0] T594;
  wire T595;
  wire T596;
  wire[4:0] T597;
  wire T598;
  wire T599;
  reg[0:0] dramBank1_valid_received_4;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[9:0] T604;
  wire T605;
  wire T606;
  wire[4:0] T607;
  wire T608;
  wire T609;
  reg[0:0] dramBank1_valid_received_3;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[9:0] T614;
  wire T615;
  wire T616;
  wire[4:0] T617;
  wire T618;
  wire T619;
  reg[0:0] dramBank1_valid_received_2;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[9:0] T624;
  wire T625;
  wire T626;
  wire[4:0] T627;
  wire T628;
  wire T629;
  reg[0:0] dramBank1_valid_received_1;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire[9:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  reg[0:0] dramBank1_valid_received_0;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire[9:0] T643;
  wire T644;
  wire T645;
  wire[4:0] T646;
  wire T647;
  wire T648;
  reg[0:0] dramBank1PortHadReadyRequest;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  reg[0:0] dramBank1_ready_received;
  wire T653;
  wire T654;
  wire dramBank1Port_req_ready;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire dramBank0Port_req_valid;
  wire T659;
  wire T660;
  wire T661;
  wire[7:0] T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  reg[0:0] dramBank0_valid_received_7;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire[9:0] T672;
  wire[9:0] dramBank0Port_rep_tag;
  wire dramBank0Port_rep_ready;
  wire[9:0] dramBank0Port_req_tag;
  wire[9:0] T673;
  wire dramBank0Port_rep_valid;
  wire T674;
  wire T675;
  wire[4:0] T676;
  wire T677;
  wire T678;
  reg[0:0] dramBank0_valid_received_6;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire[9:0] T683;
  wire T684;
  wire T685;
  wire[4:0] T686;
  wire T687;
  wire T688;
  reg[0:0] dramBank0_valid_received_5;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire[9:0] T693;
  wire T694;
  wire T695;
  wire[4:0] T696;
  wire T697;
  wire T698;
  reg[0:0] dramBank0_valid_received_4;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire[9:0] T703;
  wire T704;
  wire T705;
  wire[4:0] T706;
  wire T707;
  wire T708;
  reg[0:0] dramBank0_valid_received_3;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[9:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  reg[0:0] dramBank0_valid_received_2;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire[9:0] T723;
  wire T724;
  wire T725;
  wire[4:0] T726;
  wire T727;
  wire T728;
  reg[0:0] dramBank0_valid_received_1;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire[9:0] T733;
  wire T734;
  wire T735;
  wire[4:0] T736;
  wire T737;
  reg[0:0] dramBank0_valid_received_0;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[9:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  reg[0:0] dramBank0PortHadReadyRequest;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  reg[0:0] dramBank0_ready_received;
  wire T752;
  wire T753;
  wire dramBank0Port_req_ready;
  wire T754;
  wire T755;
  reg[0:0] subStateTh_6;
  wire T756;
  wire T757;
  wire T758;
  wire[3:0] T759;
  wire T760;
  wire T761;
  reg[7:0] State_6;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[7:0] T767;
  wire[7:0] T768;
  wire[7:0] T769;
  wire[7:0] T770;
  wire[7:0] T771;
  wire[7:0] T772;
  wire[7:0] T773;
  wire[7:0] T774;
  wire[7:0] T775;
  wire[7:0] T776;
  wire T777;
  reg[7:0] State_5;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[7:0] T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[7:0] T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[7:0] T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire[7:0] T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire[7:0] T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[7:0] T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[7:0] T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire[7:0] T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire[47:0] T833;
  wire[47:0] b;
  wire[47:0] T834;
  wire[31:0] T835;
  wire[31:0] T836;
  wire[31:0] T837;
  wire[31:0] T838;
  reg[31:0] inputReg_7_addr;
  wire T839;
  wire T840;
  wire[7:0] T841;
  wire[22:0] T842;
  wire T843;
  wire T844;
  wire[31:0] T845;
  wire[31:0] T846;
  wire[31:0] T847;
  wire[31:0] T848;
  reg[31:0] inputReg_6_addr;
  wire T849;
  wire T850;
  wire[31:0] T851;
  wire[31:0] T852;
  wire[31:0] T853;
  wire[31:0] T854;
  reg[31:0] inputReg_5_addr;
  wire T855;
  wire T856;
  wire[31:0] T857;
  wire[31:0] T858;
  wire[31:0] T859;
  wire[31:0] T860;
  wire T861;
  reg[31:0] inputReg_4_addr;
  wire T862;
  wire T863;
  wire[31:0] T864;
  wire[31:0] T865;
  wire[31:0] T866;
  wire[31:0] T867;
  wire T868;
  reg[31:0] inputReg_3_addr;
  wire T869;
  wire T870;
  wire[31:0] T871;
  wire[31:0] T872;
  wire[31:0] T873;
  wire[31:0] T874;
  wire T875;
  reg[31:0] inputReg_2_addr;
  wire T876;
  wire T877;
  wire[31:0] T878;
  wire[31:0] T879;
  wire[31:0] T880;
  wire[31:0] T881;
  wire T882;
  reg[31:0] inputReg_1_addr;
  wire T883;
  wire T884;
  wire[31:0] T885;
  wire[31:0] T886;
  wire[31:0] T887;
  wire T888;
  reg[31:0] inputReg_0_addr;
  wire T889;
  wire T890;
  wire[31:0] T891;
  wire T892;
  wire T893;
  wire T894;
  wire[47:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[47:0] T899;
  wire T900;
  wire T901;
  wire T902;
  wire[47:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[47:0] T907;
  wire T908;
  wire T909;
  wire T910;
  wire[47:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[47:0] T915;
  wire T916;
  wire T917;
  wire T918;
  wire[47:0] T919;
  wire T920;
  wire T921;
  wire[7:0] T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire T928;
  wire[59:0] r;
  wire[59:0] T929;
  wire[31:0] T930;
  wire[59:0] T931;
  wire[31:0] T932;
  wire[31:0] T933;
  wire[31:0] T934;
  reg[31:0] rb7RowAddr_7;
  wire T935;
  wire T936;
  wire[59:0] T937;
  wire[59:0] T938;
  wire[31:0] T939;
  wire[31:0] T940;
  wire[31:0] T941;
  wire[31:0] T942;
  reg[31:0] rb7RowAddr_6;
  wire T943;
  wire T944;
  wire[59:0] T945;
  wire[59:0] T946;
  wire[31:0] T947;
  wire[31:0] T948;
  wire[31:0] T949;
  wire[31:0] T950;
  reg[31:0] rb7RowAddr_5;
  wire T951;
  wire[59:0] T952;
  wire[59:0] T953;
  wire[31:0] T954;
  wire[31:0] T955;
  wire[31:0] T956;
  wire[31:0] T957;
  reg[31:0] rb7RowAddr_4;
  wire T958;
  wire T959;
  wire[59:0] T960;
  wire[59:0] T961;
  wire[31:0] T962;
  wire[31:0] T963;
  wire[31:0] T964;
  wire[31:0] T965;
  reg[31:0] rb7RowAddr_3;
  wire T966;
  wire T967;
  wire[59:0] T968;
  wire[59:0] T969;
  wire[31:0] T970;
  wire[31:0] T971;
  wire[31:0] T972;
  wire[31:0] T973;
  reg[31:0] rb7RowAddr_2;
  wire T974;
  wire T975;
  wire[59:0] T976;
  wire[59:0] T977;
  wire[31:0] T978;
  wire[31:0] T979;
  wire[31:0] T980;
  wire[31:0] T981;
  reg[31:0] rb7RowAddr_1;
  wire T982;
  wire T983;
  wire[59:0] T984;
  wire[59:0] T985;
  wire[31:0] T986;
  wire[31:0] T987;
  wire[31:0] T988;
  reg[31:0] rb7RowAddr_0;
  wire T989;
  wire T990;
  wire[59:0] T991;
  wire[59:0] T992;
  wire[31:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[59:0] T1003;
  wire[31:0] T1004;
  wire[31:0] T1005;
  wire[31:0] T1006;
  reg[31:0] rb6RowAddr_7;
  wire T1007;
  wire T1008;
  wire[59:0] T1009;
  wire[59:0] T1010;
  wire[31:0] T1011;
  wire[31:0] T1012;
  wire[31:0] T1013;
  wire[31:0] T1014;
  reg[31:0] rb6RowAddr_6;
  wire T1015;
  wire T1016;
  wire[59:0] T1017;
  wire[59:0] T1018;
  wire[31:0] T1019;
  wire[31:0] T1020;
  wire[31:0] T1021;
  wire[31:0] T1022;
  reg[31:0] rb6RowAddr_5;
  wire T1023;
  wire[59:0] T1024;
  wire[59:0] T1025;
  wire[31:0] T1026;
  wire[31:0] T1027;
  wire[31:0] T1028;
  wire[31:0] T1029;
  reg[31:0] rb6RowAddr_4;
  wire T1030;
  wire T1031;
  wire[59:0] T1032;
  wire[59:0] T1033;
  wire[31:0] T1034;
  wire[31:0] T1035;
  wire[31:0] T1036;
  wire[31:0] T1037;
  reg[31:0] rb6RowAddr_3;
  wire T1038;
  wire T1039;
  wire[59:0] T1040;
  wire[59:0] T1041;
  wire[31:0] T1042;
  wire[31:0] T1043;
  wire[31:0] T1044;
  wire[31:0] T1045;
  reg[31:0] rb6RowAddr_2;
  wire T1046;
  wire T1047;
  wire[59:0] T1048;
  wire[59:0] T1049;
  wire[31:0] T1050;
  wire[31:0] T1051;
  wire[31:0] T1052;
  wire[31:0] T1053;
  reg[31:0] rb6RowAddr_1;
  wire T1054;
  wire T1055;
  wire[59:0] T1056;
  wire[59:0] T1057;
  wire[31:0] T1058;
  wire[31:0] T1059;
  wire[31:0] T1060;
  reg[31:0] rb6RowAddr_0;
  wire T1061;
  wire T1062;
  wire[59:0] T1063;
  wire[59:0] T1064;
  wire[31:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire[59:0] T1075;
  wire[31:0] T1076;
  wire[31:0] T1077;
  wire[31:0] T1078;
  reg[31:0] rb5RowAddr_7;
  wire T1079;
  wire T1080;
  wire[59:0] T1081;
  wire[59:0] T1082;
  wire[31:0] T1083;
  wire[31:0] T1084;
  wire[31:0] T1085;
  wire[31:0] T1086;
  reg[31:0] rb5RowAddr_6;
  wire T1087;
  wire T1088;
  wire[59:0] T1089;
  wire[59:0] T1090;
  wire[31:0] T1091;
  wire[31:0] T1092;
  wire[31:0] T1093;
  wire[31:0] T1094;
  reg[31:0] rb5RowAddr_5;
  wire T1095;
  wire[59:0] T1096;
  wire[59:0] T1097;
  wire[31:0] T1098;
  wire[31:0] T1099;
  wire[31:0] T1100;
  wire[31:0] T1101;
  reg[31:0] rb5RowAddr_4;
  wire T1102;
  wire T1103;
  wire[59:0] T1104;
  wire[59:0] T1105;
  wire[31:0] T1106;
  wire[31:0] T1107;
  wire[31:0] T1108;
  wire[31:0] T1109;
  reg[31:0] rb5RowAddr_3;
  wire T1110;
  wire T1111;
  wire[59:0] T1112;
  wire[59:0] T1113;
  wire[31:0] T1114;
  wire[31:0] T1115;
  wire[31:0] T1116;
  wire[31:0] T1117;
  reg[31:0] rb5RowAddr_2;
  wire T1118;
  wire T1119;
  wire[59:0] T1120;
  wire[59:0] T1121;
  wire[31:0] T1122;
  wire[31:0] T1123;
  wire[31:0] T1124;
  wire[31:0] T1125;
  reg[31:0] rb5RowAddr_1;
  wire T1126;
  wire T1127;
  wire[59:0] T1128;
  wire[59:0] T1129;
  wire[31:0] T1130;
  wire[31:0] T1131;
  wire[31:0] T1132;
  reg[31:0] rb5RowAddr_0;
  wire T1133;
  wire T1134;
  wire[59:0] T1135;
  wire[59:0] T1136;
  wire[31:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire[59:0] T1147;
  wire[31:0] T1148;
  wire[31:0] T1149;
  wire[31:0] T1150;
  reg[31:0] rb4RowAddr_7;
  wire T1151;
  wire T1152;
  wire[59:0] T1153;
  wire[59:0] T1154;
  wire[31:0] T1155;
  wire[31:0] T1156;
  wire[31:0] T1157;
  wire[31:0] T1158;
  reg[31:0] rb4RowAddr_6;
  wire T1159;
  wire T1160;
  wire[59:0] T1161;
  wire[59:0] T1162;
  wire[31:0] T1163;
  wire[31:0] T1164;
  wire[31:0] T1165;
  wire[31:0] T1166;
  reg[31:0] rb4RowAddr_5;
  wire T1167;
  wire[59:0] T1168;
  wire[59:0] T1169;
  wire[31:0] T1170;
  wire[31:0] T1171;
  wire[31:0] T1172;
  wire[31:0] T1173;
  reg[31:0] rb4RowAddr_4;
  wire T1174;
  wire T1175;
  wire[59:0] T1176;
  wire[59:0] T1177;
  wire[31:0] T1178;
  wire[31:0] T1179;
  wire[31:0] T1180;
  wire[31:0] T1181;
  reg[31:0] rb4RowAddr_3;
  wire T1182;
  wire T1183;
  wire[59:0] T1184;
  wire[59:0] T1185;
  wire[31:0] T1186;
  wire[31:0] T1187;
  wire[31:0] T1188;
  wire[31:0] T1189;
  reg[31:0] rb4RowAddr_2;
  wire T1190;
  wire T1191;
  wire[59:0] T1192;
  wire[59:0] T1193;
  wire[31:0] T1194;
  wire[31:0] T1195;
  wire[31:0] T1196;
  wire[31:0] T1197;
  reg[31:0] rb4RowAddr_1;
  wire T1198;
  wire T1199;
  wire[59:0] T1200;
  wire[59:0] T1201;
  wire[31:0] T1202;
  wire[31:0] T1203;
  wire[31:0] T1204;
  reg[31:0] rb4RowAddr_0;
  wire T1205;
  wire T1206;
  wire[59:0] T1207;
  wire[59:0] T1208;
  wire[31:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire[59:0] T1219;
  wire[31:0] T1220;
  wire[31:0] T1221;
  wire[31:0] T1222;
  reg[31:0] rb3RowAddr_7;
  wire T1223;
  wire T1224;
  wire[59:0] T1225;
  wire[59:0] T1226;
  wire[31:0] T1227;
  wire[31:0] T1228;
  wire[31:0] T1229;
  wire[31:0] T1230;
  reg[31:0] rb3RowAddr_6;
  wire T1231;
  wire T1232;
  wire[59:0] T1233;
  wire[59:0] T1234;
  wire[31:0] T1235;
  wire[31:0] T1236;
  wire[31:0] T1237;
  wire[31:0] T1238;
  reg[31:0] rb3RowAddr_5;
  wire T1239;
  wire[59:0] T1240;
  wire[59:0] T1241;
  wire[31:0] T1242;
  wire[31:0] T1243;
  wire[31:0] T1244;
  wire[31:0] T1245;
  reg[31:0] rb3RowAddr_4;
  wire T1246;
  wire T1247;
  wire[59:0] T1248;
  wire[59:0] T1249;
  wire[31:0] T1250;
  wire[31:0] T1251;
  wire[31:0] T1252;
  wire[31:0] T1253;
  reg[31:0] rb3RowAddr_3;
  wire T1254;
  wire T1255;
  wire[59:0] T1256;
  wire[59:0] T1257;
  wire[31:0] T1258;
  wire[31:0] T1259;
  wire[31:0] T1260;
  wire[31:0] T1261;
  reg[31:0] rb3RowAddr_2;
  wire T1262;
  wire T1263;
  wire[59:0] T1264;
  wire[59:0] T1265;
  wire[31:0] T1266;
  wire[31:0] T1267;
  wire[31:0] T1268;
  wire[31:0] T1269;
  reg[31:0] rb3RowAddr_1;
  wire T1270;
  wire T1271;
  wire[59:0] T1272;
  wire[59:0] T1273;
  wire[31:0] T1274;
  wire[31:0] T1275;
  wire[31:0] T1276;
  reg[31:0] rb3RowAddr_0;
  wire T1277;
  wire T1278;
  wire[59:0] T1279;
  wire[59:0] T1280;
  wire[31:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire[59:0] T1291;
  wire[31:0] T1292;
  wire[31:0] T1293;
  wire[31:0] T1294;
  reg[31:0] rb2RowAddr_7;
  wire T1295;
  wire T1296;
  wire[59:0] T1297;
  wire[59:0] T1298;
  wire[31:0] T1299;
  wire[31:0] T1300;
  wire[31:0] T1301;
  wire[31:0] T1302;
  reg[31:0] rb2RowAddr_6;
  wire T1303;
  wire T1304;
  wire[59:0] T1305;
  wire[59:0] T1306;
  wire[31:0] T1307;
  wire[31:0] T1308;
  wire[31:0] T1309;
  wire[31:0] T1310;
  reg[31:0] rb2RowAddr_5;
  wire T1311;
  wire[59:0] T1312;
  wire[59:0] T1313;
  wire[31:0] T1314;
  wire[31:0] T1315;
  wire[31:0] T1316;
  wire[31:0] T1317;
  reg[31:0] rb2RowAddr_4;
  wire T1318;
  wire T1319;
  wire[59:0] T1320;
  wire[59:0] T1321;
  wire[31:0] T1322;
  wire[31:0] T1323;
  wire[31:0] T1324;
  wire[31:0] T1325;
  reg[31:0] rb2RowAddr_3;
  wire T1326;
  wire T1327;
  wire[59:0] T1328;
  wire[59:0] T1329;
  wire[31:0] T1330;
  wire[31:0] T1331;
  wire[31:0] T1332;
  wire[31:0] T1333;
  reg[31:0] rb2RowAddr_2;
  wire T1334;
  wire T1335;
  wire[59:0] T1336;
  wire[59:0] T1337;
  wire[31:0] T1338;
  wire[31:0] T1339;
  wire[31:0] T1340;
  wire[31:0] T1341;
  reg[31:0] rb2RowAddr_1;
  wire T1342;
  wire T1343;
  wire[59:0] T1344;
  wire[59:0] T1345;
  wire[31:0] T1346;
  wire[31:0] T1347;
  wire[31:0] T1348;
  reg[31:0] rb2RowAddr_0;
  wire T1349;
  wire T1350;
  wire[59:0] T1351;
  wire[59:0] T1352;
  wire[31:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire[59:0] T1363;
  wire[31:0] T1364;
  wire[31:0] T1365;
  wire[31:0] T1366;
  reg[31:0] rb1RowAddr_7;
  wire T1367;
  wire T1368;
  wire[59:0] T1369;
  wire[59:0] T1370;
  wire[31:0] T1371;
  wire[31:0] T1372;
  wire[31:0] T1373;
  wire[31:0] T1374;
  reg[31:0] rb1RowAddr_6;
  wire T1375;
  wire T1376;
  wire[59:0] T1377;
  wire[59:0] T1378;
  wire[31:0] T1379;
  wire[31:0] T1380;
  wire[31:0] T1381;
  wire[31:0] T1382;
  reg[31:0] rb1RowAddr_5;
  wire T1383;
  wire[59:0] T1384;
  wire[59:0] T1385;
  wire[31:0] T1386;
  wire[31:0] T1387;
  wire[31:0] T1388;
  wire[31:0] T1389;
  reg[31:0] rb1RowAddr_4;
  wire T1390;
  wire T1391;
  wire[59:0] T1392;
  wire[59:0] T1393;
  wire[31:0] T1394;
  wire[31:0] T1395;
  wire[31:0] T1396;
  wire[31:0] T1397;
  reg[31:0] rb1RowAddr_3;
  wire T1398;
  wire T1399;
  wire[59:0] T1400;
  wire[59:0] T1401;
  wire[31:0] T1402;
  wire[31:0] T1403;
  wire[31:0] T1404;
  wire[31:0] T1405;
  reg[31:0] rb1RowAddr_2;
  wire T1406;
  wire T1407;
  wire[59:0] T1408;
  wire[59:0] T1409;
  wire[31:0] T1410;
  wire[31:0] T1411;
  wire[31:0] T1412;
  wire[31:0] T1413;
  reg[31:0] rb1RowAddr_1;
  wire T1414;
  wire T1415;
  wire[59:0] T1416;
  wire[59:0] T1417;
  wire[31:0] T1418;
  wire[31:0] T1419;
  wire[31:0] T1420;
  reg[31:0] rb1RowAddr_0;
  wire T1421;
  wire T1422;
  wire[59:0] T1423;
  wire[59:0] T1424;
  wire[31:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire[59:0] T1435;
  wire[31:0] T1436;
  wire[31:0] T1437;
  wire[31:0] T1438;
  reg[31:0] rb0RowAddr_7;
  wire T1439;
  wire T1440;
  wire[59:0] T1441;
  wire[59:0] T1442;
  wire[31:0] T1443;
  wire[31:0] T1444;
  wire[31:0] T1445;
  wire[31:0] T1446;
  reg[31:0] rb0RowAddr_6;
  wire T1447;
  wire T1448;
  wire[59:0] T1449;
  wire[59:0] T1450;
  wire[31:0] T1451;
  wire[31:0] T1452;
  wire[31:0] T1453;
  wire[31:0] T1454;
  reg[31:0] rb0RowAddr_5;
  wire T1455;
  wire[59:0] T1456;
  wire[59:0] T1457;
  wire[31:0] T1458;
  wire[31:0] T1459;
  wire[31:0] T1460;
  wire[31:0] T1461;
  reg[31:0] rb0RowAddr_4;
  wire T1462;
  wire T1463;
  wire[59:0] T1464;
  wire[59:0] T1465;
  wire[31:0] T1466;
  wire[31:0] T1467;
  wire[31:0] T1468;
  wire[31:0] T1469;
  reg[31:0] rb0RowAddr_3;
  wire T1470;
  wire T1471;
  wire[59:0] T1472;
  wire[59:0] T1473;
  wire[31:0] T1474;
  wire[31:0] T1475;
  wire[31:0] T1476;
  wire[31:0] T1477;
  reg[31:0] rb0RowAddr_2;
  wire T1478;
  wire T1479;
  wire[59:0] T1480;
  wire[59:0] T1481;
  wire[31:0] T1482;
  wire[31:0] T1483;
  wire[31:0] T1484;
  wire[31:0] T1485;
  reg[31:0] rb0RowAddr_1;
  wire T1486;
  wire T1487;
  wire[59:0] T1488;
  wire[59:0] T1489;
  wire[31:0] T1490;
  wire[31:0] T1491;
  wire[31:0] T1492;
  reg[31:0] rb0RowAddr_0;
  wire T1493;
  wire T1494;
  wire[59:0] T1495;
  wire[59:0] T1496;
  wire[31:0] T1497;
  wire T1498;
  wire T1499;
  wire T1500;
  wire T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire[7:0] T1508;
  wire[7:0] T1509;
  wire[7:0] T1510;
  wire[7:0] T1511;
  wire[7:0] T1512;
  wire[7:0] T1513;
  wire[7:0] T1514;
  wire[7:0] T1515;
  wire[7:0] T1516;
  wire[7:0] T1517;
  wire[7:0] T1518;
  wire[7:0] T1519;
  wire[7:0] T1520;
  wire[7:0] T1521;
  wire[7:0] T1522;
  wire[7:0] T1523;
  wire[7:0] T1524;
  wire[7:0] T1525;
  wire[7:0] T1526;
  wire[7:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[7:0] T1530;
  wire[7:0] T1531;
  reg[7:0] EmitReturnState_7;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  wire T1546;
  wire T1547;
  wire[7:0] T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire T1556;
  wire[7:0] T1557;
  wire[7:0] T1558;
  wire[7:0] T1559;
  reg[7:0] EmitReturnState_6;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire[7:0] T1576;
  wire T1577;
  wire T1578;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[7:0] T1585;
  wire[7:0] T1586;
  wire[7:0] T1587;
  reg[7:0] EmitReturnState_5;
  wire T1588;
  wire T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire[7:0] T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire T1604;
  wire[7:0] T1605;
  wire[7:0] T1606;
  wire[7:0] T1607;
  reg[7:0] EmitReturnState_4;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire T1620;
  wire T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[7:0] T1625;
  wire T1626;
  wire T1627;
  wire T1628;
  wire T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire[7:0] T1634;
  wire[7:0] T1635;
  wire[7:0] T1636;
  reg[7:0] EmitReturnState_3;
  wire T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire T1644;
  wire T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire T1652;
  wire T1653;
  wire[7:0] T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire[7:0] T1663;
  wire[7:0] T1664;
  wire[7:0] T1665;
  reg[7:0] EmitReturnState_2;
  wire T1666;
  wire T1667;
  wire T1668;
  wire T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire T1676;
  wire T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire[7:0] T1683;
  wire T1684;
  wire T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire T1689;
  wire T1690;
  wire T1691;
  wire[7:0] T1692;
  wire[7:0] T1693;
  wire[7:0] T1694;
  reg[7:0] EmitReturnState_1;
  wire T1695;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire T1700;
  wire T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire T1705;
  wire T1706;
  wire T1707;
  wire T1708;
  wire T1709;
  wire T1710;
  wire T1711;
  wire[7:0] T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire T1716;
  wire T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[7:0] T1721;
  wire[7:0] T1722;
  reg[7:0] EmitReturnState_0;
  wire T1723;
  wire T1724;
  wire T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire T1738;
  wire T1739;
  wire[7:0] T1740;
  wire T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire T1745;
  wire T1746;
  wire T1747;
  wire T1748;
  wire[7:0] T1749;
  wire[7:0] T1750;
  wire[7:0] T1751;
  wire[7:0] T1752;
  wire[7:0] T1753;
  wire[7:0] T1754;
  wire[7:0] T1755;
  wire[7:0] T1756;
  wire[7:0] T1757;
  wire[7:0] T1758;
  wire[7:0] T1759;
  wire[7:0] T1760;
  wire[7:0] T1761;
  wire[7:0] T1762;
  wire[7:0] T1763;
  wire[7:0] T1764;
  wire[7:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire T1770;
  wire T1771;
  wire T1772;
  wire T1773;
  wire[7:0] T1774;
  wire[7:0] T1775;
  wire[7:0] T1776;
  reg[7:0] State_4;
  wire T1777;
  wire T1778;
  wire T1779;
  wire T1780;
  wire T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire T1788;
  wire T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire T1796;
  wire T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire T1804;
  wire T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire T1812;
  wire T1813;
  wire[7:0] T1814;
  wire[7:0] T1815;
  wire[7:0] T1816;
  wire[7:0] T1817;
  wire[7:0] T1818;
  wire[7:0] T1819;
  wire[7:0] T1820;
  wire[7:0] T1821;
  wire[7:0] T1822;
  wire[7:0] T1823;
  wire[7:0] T1824;
  wire[7:0] T1825;
  wire[7:0] T1826;
  wire[7:0] T1827;
  wire[7:0] T1828;
  wire[7:0] T1829;
  wire[7:0] T1830;
  wire[7:0] T1831;
  wire[7:0] T1832;
  wire[7:0] T1833;
  wire[7:0] T1834;
  wire[7:0] T1835;
  wire[7:0] T1836;
  wire[7:0] T1837;
  wire[7:0] T1838;
  wire[7:0] T1839;
  wire[7:0] T1840;
  wire[7:0] T1841;
  wire[7:0] T1842;
  wire[7:0] T1843;
  wire[7:0] T1844;
  wire[7:0] T1845;
  wire[7:0] T1846;
  wire[7:0] T1847;
  wire[7:0] T1848;
  wire[7:0] T1849;
  wire[7:0] T1850;
  wire[7:0] T1851;
  wire T1852;
  wire T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire T1859;
  wire[7:0] T1860;
  wire[7:0] T1861;
  wire[7:0] T1862;
  reg[7:0] State_3;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire T1868;
  wire T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire T1884;
  wire T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[7:0] T1900;
  wire[7:0] T1901;
  wire[7:0] T1902;
  wire[7:0] T1903;
  wire[7:0] T1904;
  wire[7:0] T1905;
  wire[7:0] T1906;
  wire[7:0] T1907;
  wire[7:0] T1908;
  wire[7:0] T1909;
  wire[7:0] T1910;
  wire[7:0] T1911;
  wire[7:0] T1912;
  wire[7:0] T1913;
  wire[7:0] T1914;
  wire[7:0] T1915;
  wire[7:0] T1916;
  wire[7:0] T1917;
  wire[7:0] T1918;
  wire[7:0] T1919;
  wire[7:0] T1920;
  wire[7:0] T1921;
  wire[7:0] T1922;
  wire[7:0] T1923;
  wire[7:0] T1924;
  wire[7:0] T1925;
  wire[7:0] T1926;
  wire[7:0] T1927;
  wire[7:0] T1928;
  wire[7:0] T1929;
  wire[7:0] T1930;
  wire[7:0] T1931;
  wire[7:0] T1932;
  wire[7:0] T1933;
  wire[7:0] T1934;
  wire[7:0] T1935;
  wire[7:0] T1936;
  wire[7:0] T1937;
  wire T1938;
  wire T1939;
  wire T1940;
  wire T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire T1945;
  wire[7:0] T1946;
  wire[7:0] T1947;
  wire[7:0] T1948;
  reg[7:0] State_2;
  wire T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire T1955;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  wire T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire T1985;
  wire[7:0] T1986;
  wire[7:0] T1987;
  wire[7:0] T1988;
  wire[7:0] T1989;
  wire[7:0] T1990;
  wire[7:0] T1991;
  wire[7:0] T1992;
  wire[7:0] T1993;
  wire[7:0] T1994;
  wire[7:0] T1995;
  wire[7:0] T1996;
  wire[7:0] T1997;
  wire[7:0] T1998;
  wire[7:0] T1999;
  wire[7:0] T2000;
  wire[7:0] T2001;
  wire[7:0] T2002;
  wire[7:0] T2003;
  wire[7:0] T2004;
  wire[7:0] T2005;
  wire[7:0] T2006;
  wire[7:0] T2007;
  wire[7:0] T2008;
  wire[7:0] T2009;
  wire[7:0] T2010;
  wire[7:0] T2011;
  wire[7:0] T2012;
  wire[7:0] T2013;
  wire[7:0] T2014;
  wire[7:0] T2015;
  wire[7:0] T2016;
  wire[7:0] T2017;
  wire[7:0] T2018;
  wire[7:0] T2019;
  wire[7:0] T2020;
  wire[7:0] T2021;
  wire[7:0] T2022;
  wire[7:0] T2023;
  wire T2024;
  wire T2025;
  wire T2026;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire[7:0] T2032;
  wire[7:0] T2033;
  wire[7:0] T2034;
  reg[7:0] State_1;
  wire T2035;
  wire T2036;
  wire T2037;
  wire T2038;
  wire T2039;
  wire T2040;
  wire T2041;
  wire T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  wire T2051;
  wire T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  wire T2057;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire T2065;
  wire T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire T2070;
  wire T2071;
  wire[7:0] T2072;
  wire[7:0] T2073;
  wire[7:0] T2074;
  wire[7:0] T2075;
  wire[7:0] T2076;
  wire[7:0] T2077;
  wire[7:0] T2078;
  wire[7:0] T2079;
  wire[7:0] T2080;
  wire[7:0] T2081;
  wire[7:0] T2082;
  wire[7:0] T2083;
  wire[7:0] T2084;
  wire[7:0] T2085;
  wire[7:0] T2086;
  wire[7:0] T2087;
  wire[7:0] T2088;
  wire[7:0] T2089;
  wire[7:0] T2090;
  wire[7:0] T2091;
  wire[7:0] T2092;
  wire[7:0] T2093;
  wire[7:0] T2094;
  wire[7:0] T2095;
  wire[7:0] T2096;
  wire[7:0] T2097;
  wire[7:0] T2098;
  wire[7:0] T2099;
  wire[7:0] T2100;
  wire[7:0] T2101;
  wire[7:0] T2102;
  wire[7:0] T2103;
  wire[7:0] T2104;
  wire[7:0] T2105;
  wire[7:0] T2106;
  wire[7:0] T2107;
  wire[7:0] T2108;
  wire[7:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire T2116;
  wire T2117;
  wire[7:0] T2118;
  wire[7:0] T2119;
  reg[7:0] State_0;
  wire T2120;
  wire T2121;
  wire T2122;
  wire T2123;
  wire T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire T2139;
  wire T2140;
  wire T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire[7:0] T2157;
  wire[7:0] T2158;
  wire[7:0] T2159;
  wire[7:0] T2160;
  wire[7:0] T2161;
  wire[7:0] T2162;
  wire[7:0] T2163;
  wire[7:0] T2164;
  wire[7:0] T2165;
  wire[7:0] T2166;
  wire[7:0] T2167;
  wire[7:0] T2168;
  wire[7:0] T2169;
  wire[7:0] T2170;
  wire[7:0] T2171;
  wire[7:0] T2172;
  wire[7:0] T2173;
  wire[7:0] T2174;
  wire[7:0] T2175;
  wire[7:0] T2176;
  wire[7:0] T2177;
  wire[7:0] T2178;
  wire[7:0] T2179;
  wire[7:0] T2180;
  wire[7:0] T2181;
  wire[7:0] T2182;
  wire[7:0] T2183;
  wire[7:0] T2184;
  wire[7:0] T2185;
  wire[7:0] T2186;
  wire[7:0] T2187;
  wire[7:0] T2188;
  wire[7:0] T2189;
  wire[7:0] T2190;
  wire[7:0] T2191;
  wire[7:0] T2192;
  wire[7:0] T2193;
  wire[7:0] T2194;
  wire T2195;
  wire T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire T2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  wire T2211;
  wire T2212;
  wire T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire T2225;
  wire T2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  wire T2236;
  wire T2237;
  wire T2238;
  wire T2239;
  wire[7:0] T2240;
  wire[7:0] T2241;
  wire[7:0] T2242;
  wire[7:0] T2243;
  wire[7:0] T2244;
  wire[7:0] T2245;
  wire[7:0] T2246;
  wire[7:0] T2247;
  wire[7:0] T2248;
  wire[7:0] T2249;
  wire[7:0] T2250;
  wire[7:0] T2251;
  wire[7:0] T2252;
  wire[7:0] T2253;
  wire[7:0] T2254;
  wire[7:0] T2255;
  wire[7:0] T2256;
  wire[7:0] T2257;
  wire[7:0] T2258;
  wire[7:0] T2259;
  wire[7:0] T2260;
  wire[7:0] T2261;
  wire[7:0] T2262;
  wire[7:0] T2263;
  wire[7:0] T2264;
  wire[7:0] T2265;
  wire[7:0] T2266;
  wire[7:0] T2267;
  wire[7:0] T2268;
  wire[7:0] T2269;
  wire[7:0] T2270;
  wire[7:0] T2271;
  wire[7:0] T2272;
  wire[7:0] T2273;
  wire[7:0] T2274;
  wire[7:0] T2275;
  wire[7:0] T2276;
  wire[7:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire T2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire T2289;
  wire[3:0] T2290;
  wire T2291;
  reg[0:0] subStateTh_5;
  wire T2292;
  wire T2293;
  wire T2294;
  wire[3:0] T2295;
  wire T2296;
  wire T2297;
  wire T2298;
  wire T2299;
  wire T2300;
  wire T2301;
  wire[3:0] T2302;
  wire T2303;
  reg[0:0] subStateTh_4;
  wire T2304;
  wire T2305;
  wire T2306;
  wire[3:0] T2307;
  wire T2308;
  wire T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire T2313;
  wire[3:0] T2314;
  wire T2315;
  reg[0:0] subStateTh_3;
  wire T2316;
  wire T2317;
  wire T2318;
  wire[3:0] T2319;
  wire T2320;
  wire T2321;
  wire T2322;
  wire T2323;
  wire T2324;
  wire T2325;
  wire[3:0] T2326;
  wire T2327;
  reg[0:0] subStateTh_2;
  wire T2328;
  wire T2329;
  wire T2330;
  wire[3:0] T2331;
  wire T2332;
  wire T2333;
  wire T2334;
  wire T2335;
  wire T2336;
  wire T2337;
  wire[3:0] T2338;
  wire T2339;
  reg[0:0] subStateTh_1;
  wire T2340;
  wire T2341;
  wire T2342;
  wire[3:0] T2343;
  wire T2344;
  wire T2345;
  wire T2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire[3:0] T2350;
  wire T2351;
  reg[0:0] subStateTh_0;
  wire T2352;
  wire T2353;
  wire T2354;
  wire[3:0] T2355;
  wire T2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  wire T2361;
  wire[3:0] T2362;
  wire T2363;
  wire[7:0] T2364;
  wire[7:0] T2365;
  wire[7:0] T2366;
  wire[7:0] T2367;
  wire[7:0] T2368;
  wire[7:0] T2369;
  wire[7:0] T2370;
  wire[7:0] T2371;
  wire[7:0] T2372;
  wire[7:0] T2373;
  wire[7:0] T2374;
  wire[7:0] T2375;
  wire[7:0] T2376;
  wire[7:0] T2377;
  wire[7:0] T2378;
  wire[7:0] T2379;
  wire[7:0] T2380;
  wire[7:0] T2381;
  wire[7:0] T2382;
  wire[7:0] T2383;
  wire T2384;
  wire T2385;
  wire T2386;
  wire T2387;
  wire T2388;
  reg[0:0] dramBank7_valid_received_7;
  wire T2389;
  wire T2390;
  wire T2391;
  wire T2392;
  wire[9:0] T2393;
  wire[9:0] dramBank7Port_rep_tag;
  wire[9:0] dramBank7Port_req_tag;
  wire[9:0] T2394;
  wire dramBank7Port_rep_valid;
  wire T2395;
  wire T2396;
  wire[4:0] T2397;
  wire T2398;
  wire T2399;
  reg[0:0] dramBank7_valid_received_6;
  wire T2400;
  wire T2401;
  wire T2402;
  wire T2403;
  wire[9:0] T2404;
  wire T2405;
  wire T2406;
  wire[4:0] T2407;
  wire T2408;
  wire T2409;
  reg[0:0] dramBank7_valid_received_5;
  wire T2410;
  wire T2411;
  wire T2412;
  wire T2413;
  wire[9:0] T2414;
  wire T2415;
  wire T2416;
  wire[4:0] T2417;
  wire T2418;
  wire T2419;
  reg[0:0] dramBank7_valid_received_4;
  wire T2420;
  wire T2421;
  wire T2422;
  wire T2423;
  wire[9:0] T2424;
  wire T2425;
  wire T2426;
  wire[4:0] T2427;
  wire T2428;
  wire T2429;
  reg[0:0] dramBank7_valid_received_3;
  wire T2430;
  wire T2431;
  wire T2432;
  wire T2433;
  wire[9:0] T2434;
  wire T2435;
  wire T2436;
  wire[4:0] T2437;
  wire T2438;
  wire T2439;
  reg[0:0] dramBank7_valid_received_2;
  wire T2440;
  wire T2441;
  wire T2442;
  wire T2443;
  wire[9:0] T2444;
  wire T2445;
  wire T2446;
  wire[4:0] T2447;
  wire T2448;
  wire T2449;
  reg[0:0] dramBank7_valid_received_1;
  wire T2450;
  wire T2451;
  wire T2452;
  wire T2453;
  wire[9:0] T2454;
  wire T2455;
  wire T2456;
  wire[4:0] T2457;
  wire T2458;
  reg[0:0] dramBank7_valid_received_0;
  wire T2459;
  wire T2460;
  wire T2461;
  wire T2462;
  wire[9:0] T2463;
  wire T2464;
  wire T2465;
  wire[4:0] T2466;
  wire T2467;
  wire T2468;
  wire[4:0] T2469;
  wire T2470;
  wire T2471;
  wire[4:0] T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  wire[9:0] T2476;
  wire T2477;
  wire T2478;
  wire T2479;
  reg[0:0] dramBank6PortHadValidRequest_7;
  wire T2480;
  wire T2481;
  wire T2482;
  wire T2483;
  wire[4:0] T2484;
  wire T2485;
  wire T2486;
  wire[4:0] T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  wire[9:0] T2491;
  wire T2492;
  wire T2493;
  wire T2494;
  reg[0:0] dramBank5PortHadValidRequest_7;
  wire T2495;
  wire T2496;
  wire T2497;
  wire T2498;
  wire[4:0] T2499;
  wire T2500;
  wire T2501;
  wire[4:0] T2502;
  wire T2503;
  wire T2504;
  wire T2505;
  wire[9:0] T2506;
  wire T2507;
  wire T2508;
  wire T2509;
  reg[0:0] dramBank4PortHadValidRequest_7;
  wire T2510;
  wire T2511;
  wire T2512;
  wire T2513;
  wire[4:0] T2514;
  wire T2515;
  wire T2516;
  wire[4:0] T2517;
  wire T2518;
  wire T2519;
  wire T2520;
  wire[9:0] T2521;
  wire T2522;
  wire T2523;
  wire T2524;
  reg[0:0] dramBank3PortHadValidRequest_7;
  wire T2525;
  wire T2526;
  wire T2527;
  wire T2528;
  wire[4:0] T2529;
  wire T2530;
  wire T2531;
  wire[4:0] T2532;
  wire T2533;
  wire T2534;
  wire T2535;
  wire[9:0] T2536;
  wire T2537;
  wire T2538;
  wire T2539;
  reg[0:0] dramBank2PortHadValidRequest_7;
  wire T2540;
  wire T2541;
  wire T2542;
  wire T2543;
  wire[4:0] T2544;
  wire T2545;
  wire T2546;
  wire[4:0] T2547;
  wire T2548;
  wire T2549;
  wire T2550;
  wire[9:0] T2551;
  wire T2552;
  wire T2553;
  wire T2554;
  reg[0:0] dramBank1PortHadValidRequest_7;
  wire T2555;
  wire T2556;
  wire T2557;
  wire T2558;
  wire[4:0] T2559;
  wire T2560;
  wire T2561;
  wire[4:0] T2562;
  wire T2563;
  wire T2564;
  wire T2565;
  wire[9:0] T2566;
  wire T2567;
  wire T2568;
  reg[0:0] dramBank0PortHadValidRequest_7;
  wire T2569;
  wire T2570;
  wire T2571;
  wire T2572;
  wire[4:0] T2573;
  wire T2574;
  wire T2575;
  wire[4:0] T2576;
  wire T2577;
  wire T2578;
  wire T2579;
  wire[9:0] T2580;
  wire T2581;
  wire T2582;
  wire AllOffloadsValid_6;
  wire T2583;
  wire T2584;
  wire T2585;
  reg[0:0] dramBank7PortHadValidRequest_6;
  wire T2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire[4:0] T2590;
  wire T2591;
  wire T2592;
  wire[4:0] T2593;
  wire T2594;
  wire T2595;
  wire T2596;
  wire[9:0] T2597;
  wire T2598;
  wire T2599;
  wire T2600;
  reg[0:0] dramBank6PortHadValidRequest_6;
  wire T2601;
  wire T2602;
  wire T2603;
  wire T2604;
  wire[4:0] T2605;
  wire T2606;
  wire T2607;
  wire[4:0] T2608;
  wire T2609;
  wire T2610;
  wire T2611;
  wire[9:0] T2612;
  wire T2613;
  wire T2614;
  wire T2615;
  reg[0:0] dramBank5PortHadValidRequest_6;
  wire T2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire[4:0] T2620;
  wire T2621;
  wire T2622;
  wire[4:0] T2623;
  wire T2624;
  wire T2625;
  wire T2626;
  wire[9:0] T2627;
  wire T2628;
  wire T2629;
  wire T2630;
  reg[0:0] dramBank4PortHadValidRequest_6;
  wire T2631;
  wire T2632;
  wire T2633;
  wire T2634;
  wire[4:0] T2635;
  wire T2636;
  wire T2637;
  wire[4:0] T2638;
  wire T2639;
  wire T2640;
  wire T2641;
  wire[9:0] T2642;
  wire T2643;
  wire T2644;
  wire T2645;
  reg[0:0] dramBank3PortHadValidRequest_6;
  wire T2646;
  wire T2647;
  wire T2648;
  wire T2649;
  wire[4:0] T2650;
  wire T2651;
  wire T2652;
  wire[4:0] T2653;
  wire T2654;
  wire T2655;
  wire T2656;
  wire[9:0] T2657;
  wire T2658;
  wire T2659;
  wire T2660;
  reg[0:0] dramBank2PortHadValidRequest_6;
  wire T2661;
  wire T2662;
  wire T2663;
  wire T2664;
  wire[4:0] T2665;
  wire T2666;
  wire T2667;
  wire[4:0] T2668;
  wire T2669;
  wire T2670;
  wire T2671;
  wire[9:0] T2672;
  wire T2673;
  wire T2674;
  wire T2675;
  reg[0:0] dramBank1PortHadValidRequest_6;
  wire T2676;
  wire T2677;
  wire T2678;
  wire T2679;
  wire[4:0] T2680;
  wire T2681;
  wire T2682;
  wire[4:0] T2683;
  wire T2684;
  wire T2685;
  wire T2686;
  wire[9:0] T2687;
  wire T2688;
  wire T2689;
  reg[0:0] dramBank0PortHadValidRequest_6;
  wire T2690;
  wire T2691;
  wire T2692;
  wire T2693;
  wire[4:0] T2694;
  wire T2695;
  wire T2696;
  wire[4:0] T2697;
  wire T2698;
  wire T2699;
  wire T2700;
  wire[9:0] T2701;
  wire T2702;
  wire T2703;
  wire AllOffloadsValid_5;
  wire T2704;
  wire T2705;
  wire T2706;
  reg[0:0] dramBank7PortHadValidRequest_5;
  wire T2707;
  wire T2708;
  wire T2709;
  wire T2710;
  wire[4:0] T2711;
  wire T2712;
  wire T2713;
  wire[4:0] T2714;
  wire T2715;
  wire T2716;
  wire T2717;
  wire[9:0] T2718;
  wire T2719;
  wire T2720;
  wire T2721;
  reg[0:0] dramBank6PortHadValidRequest_5;
  wire T2722;
  wire T2723;
  wire T2724;
  wire T2725;
  wire[4:0] T2726;
  wire T2727;
  wire T2728;
  wire[4:0] T2729;
  wire T2730;
  wire T2731;
  wire T2732;
  wire[9:0] T2733;
  wire T2734;
  wire T2735;
  wire T2736;
  reg[0:0] dramBank5PortHadValidRequest_5;
  wire T2737;
  wire T2738;
  wire T2739;
  wire T2740;
  wire[4:0] T2741;
  wire T2742;
  wire T2743;
  wire[4:0] T2744;
  wire T2745;
  wire T2746;
  wire T2747;
  wire[9:0] T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  reg[0:0] dramBank4PortHadValidRequest_5;
  wire T2752;
  wire T2753;
  wire T2754;
  wire T2755;
  wire[4:0] T2756;
  wire T2757;
  wire T2758;
  wire[4:0] T2759;
  wire T2760;
  wire T2761;
  wire T2762;
  wire[9:0] T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  reg[0:0] dramBank3PortHadValidRequest_5;
  wire T2767;
  wire T2768;
  wire T2769;
  wire T2770;
  wire[4:0] T2771;
  wire T2772;
  wire T2773;
  wire[4:0] T2774;
  wire T2775;
  wire T2776;
  wire T2777;
  wire[9:0] T2778;
  wire T2779;
  wire T2780;
  wire T2781;
  reg[0:0] dramBank2PortHadValidRequest_5;
  wire T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  wire[4:0] T2786;
  wire T2787;
  wire T2788;
  wire[4:0] T2789;
  wire T2790;
  wire T2791;
  wire T2792;
  wire[9:0] T2793;
  wire T2794;
  wire T2795;
  wire T2796;
  reg[0:0] dramBank1PortHadValidRequest_5;
  wire T2797;
  wire T2798;
  wire T2799;
  wire T2800;
  wire[4:0] T2801;
  wire T2802;
  wire T2803;
  wire[4:0] T2804;
  wire T2805;
  wire T2806;
  wire T2807;
  wire[9:0] T2808;
  wire T2809;
  wire T2810;
  reg[0:0] dramBank0PortHadValidRequest_5;
  wire T2811;
  wire T2812;
  wire T2813;
  wire T2814;
  wire[4:0] T2815;
  wire T2816;
  wire T2817;
  wire[4:0] T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire[9:0] T2822;
  wire T2823;
  wire T2824;
  wire AllOffloadsValid_4;
  wire T2825;
  wire T2826;
  wire T2827;
  reg[0:0] dramBank7PortHadValidRequest_4;
  wire T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire[4:0] T2832;
  wire T2833;
  wire T2834;
  wire[4:0] T2835;
  wire T2836;
  wire T2837;
  wire T2838;
  wire[9:0] T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  reg[0:0] dramBank6PortHadValidRequest_4;
  wire T2843;
  wire T2844;
  wire T2845;
  wire T2846;
  wire[4:0] T2847;
  wire T2848;
  wire T2849;
  wire[4:0] T2850;
  wire T2851;
  wire T2852;
  wire T2853;
  wire[9:0] T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  reg[0:0] dramBank5PortHadValidRequest_4;
  wire T2858;
  wire T2859;
  wire T2860;
  wire T2861;
  wire[4:0] T2862;
  wire T2863;
  wire T2864;
  wire[4:0] T2865;
  wire T2866;
  wire T2867;
  wire T2868;
  wire[9:0] T2869;
  wire T2870;
  wire T2871;
  wire T2872;
  reg[0:0] dramBank4PortHadValidRequest_4;
  wire T2873;
  wire T2874;
  wire T2875;
  wire T2876;
  wire[4:0] T2877;
  wire T2878;
  wire T2879;
  wire[4:0] T2880;
  wire T2881;
  wire T2882;
  wire T2883;
  wire[9:0] T2884;
  wire T2885;
  wire T2886;
  wire T2887;
  reg[0:0] dramBank3PortHadValidRequest_4;
  wire T2888;
  wire T2889;
  wire T2890;
  wire T2891;
  wire[4:0] T2892;
  wire T2893;
  wire T2894;
  wire[4:0] T2895;
  wire T2896;
  wire T2897;
  wire T2898;
  wire[9:0] T2899;
  wire T2900;
  wire T2901;
  wire T2902;
  reg[0:0] dramBank2PortHadValidRequest_4;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire[4:0] T2907;
  wire T2908;
  wire T2909;
  wire[4:0] T2910;
  wire T2911;
  wire T2912;
  wire T2913;
  wire[9:0] T2914;
  wire T2915;
  wire T2916;
  wire T2917;
  reg[0:0] dramBank1PortHadValidRequest_4;
  wire T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire[4:0] T2922;
  wire T2923;
  wire T2924;
  wire[4:0] T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire[9:0] T2929;
  wire T2930;
  wire T2931;
  reg[0:0] dramBank0PortHadValidRequest_4;
  wire T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire[4:0] T2936;
  wire T2937;
  wire T2938;
  wire[4:0] T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire[9:0] T2943;
  wire T2944;
  wire T2945;
  wire AllOffloadsValid_3;
  wire T2946;
  wire T2947;
  wire T2948;
  reg[0:0] dramBank7PortHadValidRequest_3;
  wire T2949;
  wire T2950;
  wire T2951;
  wire T2952;
  wire[4:0] T2953;
  wire T2954;
  wire T2955;
  wire[4:0] T2956;
  wire T2957;
  wire T2958;
  wire T2959;
  wire[9:0] T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  reg[0:0] dramBank6PortHadValidRequest_3;
  wire T2964;
  wire T2965;
  wire T2966;
  wire T2967;
  wire[4:0] T2968;
  wire T2969;
  wire T2970;
  wire[4:0] T2971;
  wire T2972;
  wire T2973;
  wire T2974;
  wire[9:0] T2975;
  wire T2976;
  wire T2977;
  wire T2978;
  reg[0:0] dramBank5PortHadValidRequest_3;
  wire T2979;
  wire T2980;
  wire T2981;
  wire T2982;
  wire[4:0] T2983;
  wire T2984;
  wire T2985;
  wire[4:0] T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire[9:0] T2990;
  wire T2991;
  wire T2992;
  wire T2993;
  reg[0:0] dramBank4PortHadValidRequest_3;
  wire T2994;
  wire T2995;
  wire T2996;
  wire T2997;
  wire[4:0] T2998;
  wire T2999;
  wire T3000;
  wire[4:0] T3001;
  wire T3002;
  wire T3003;
  wire T3004;
  wire[9:0] T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  reg[0:0] dramBank3PortHadValidRequest_3;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire[4:0] T3013;
  wire T3014;
  wire T3015;
  wire[4:0] T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire[9:0] T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  reg[0:0] dramBank2PortHadValidRequest_3;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire[4:0] T3028;
  wire T3029;
  wire T3030;
  wire[4:0] T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire[9:0] T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  reg[0:0] dramBank1PortHadValidRequest_3;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire[4:0] T3043;
  wire T3044;
  wire T3045;
  wire[4:0] T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire[9:0] T3050;
  wire T3051;
  wire T3052;
  reg[0:0] dramBank0PortHadValidRequest_3;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire[4:0] T3057;
  wire T3058;
  wire T3059;
  wire[4:0] T3060;
  wire T3061;
  wire T3062;
  wire T3063;
  wire[9:0] T3064;
  wire T3065;
  wire T3066;
  wire AllOffloadsValid_2;
  wire T3067;
  wire T3068;
  wire T3069;
  reg[0:0] dramBank7PortHadValidRequest_2;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire[4:0] T3074;
  wire T3075;
  wire T3076;
  wire[4:0] T3077;
  wire T3078;
  wire T3079;
  wire T3080;
  wire[9:0] T3081;
  wire T3082;
  wire T3083;
  wire T3084;
  reg[0:0] dramBank6PortHadValidRequest_2;
  wire T3085;
  wire T3086;
  wire T3087;
  wire T3088;
  wire[4:0] T3089;
  wire T3090;
  wire T3091;
  wire[4:0] T3092;
  wire T3093;
  wire T3094;
  wire T3095;
  wire[9:0] T3096;
  wire T3097;
  wire T3098;
  wire T3099;
  reg[0:0] dramBank5PortHadValidRequest_2;
  wire T3100;
  wire T3101;
  wire T3102;
  wire T3103;
  wire[4:0] T3104;
  wire T3105;
  wire T3106;
  wire[4:0] T3107;
  wire T3108;
  wire T3109;
  wire T3110;
  wire[9:0] T3111;
  wire T3112;
  wire T3113;
  wire T3114;
  reg[0:0] dramBank4PortHadValidRequest_2;
  wire T3115;
  wire T3116;
  wire T3117;
  wire T3118;
  wire[4:0] T3119;
  wire T3120;
  wire T3121;
  wire[4:0] T3122;
  wire T3123;
  wire T3124;
  wire T3125;
  wire[9:0] T3126;
  wire T3127;
  wire T3128;
  wire T3129;
  reg[0:0] dramBank3PortHadValidRequest_2;
  wire T3130;
  wire T3131;
  wire T3132;
  wire T3133;
  wire[4:0] T3134;
  wire T3135;
  wire T3136;
  wire[4:0] T3137;
  wire T3138;
  wire T3139;
  wire T3140;
  wire[9:0] T3141;
  wire T3142;
  wire T3143;
  wire T3144;
  reg[0:0] dramBank2PortHadValidRequest_2;
  wire T3145;
  wire T3146;
  wire T3147;
  wire T3148;
  wire[4:0] T3149;
  wire T3150;
  wire T3151;
  wire[4:0] T3152;
  wire T3153;
  wire T3154;
  wire T3155;
  wire[9:0] T3156;
  wire T3157;
  wire T3158;
  wire T3159;
  reg[0:0] dramBank1PortHadValidRequest_2;
  wire T3160;
  wire T3161;
  wire T3162;
  wire T3163;
  wire[4:0] T3164;
  wire T3165;
  wire T3166;
  wire[4:0] T3167;
  wire T3168;
  wire T3169;
  wire T3170;
  wire[9:0] T3171;
  wire T3172;
  wire T3173;
  reg[0:0] dramBank0PortHadValidRequest_2;
  wire T3174;
  wire T3175;
  wire T3176;
  wire T3177;
  wire[4:0] T3178;
  wire T3179;
  wire T3180;
  wire[4:0] T3181;
  wire T3182;
  wire T3183;
  wire T3184;
  wire[9:0] T3185;
  wire T3186;
  wire T3187;
  wire AllOffloadsValid_1;
  wire T3188;
  wire T3189;
  wire T3190;
  reg[0:0] dramBank7PortHadValidRequest_1;
  wire T3191;
  wire T3192;
  wire T3193;
  wire T3194;
  wire[4:0] T3195;
  wire T3196;
  wire T3197;
  wire[4:0] T3198;
  wire T3199;
  wire T3200;
  wire T3201;
  wire[9:0] T3202;
  wire T3203;
  wire T3204;
  wire T3205;
  reg[0:0] dramBank6PortHadValidRequest_1;
  wire T3206;
  wire T3207;
  wire T3208;
  wire T3209;
  wire[4:0] T3210;
  wire T3211;
  wire T3212;
  wire[4:0] T3213;
  wire T3214;
  wire T3215;
  wire T3216;
  wire[9:0] T3217;
  wire T3218;
  wire T3219;
  wire T3220;
  reg[0:0] dramBank5PortHadValidRequest_1;
  wire T3221;
  wire T3222;
  wire T3223;
  wire T3224;
  wire[4:0] T3225;
  wire T3226;
  wire T3227;
  wire[4:0] T3228;
  wire T3229;
  wire T3230;
  wire T3231;
  wire[9:0] T3232;
  wire T3233;
  wire T3234;
  wire T3235;
  reg[0:0] dramBank4PortHadValidRequest_1;
  wire T3236;
  wire T3237;
  wire T3238;
  wire T3239;
  wire[4:0] T3240;
  wire T3241;
  wire T3242;
  wire[4:0] T3243;
  wire T3244;
  wire T3245;
  wire T3246;
  wire[9:0] T3247;
  wire T3248;
  wire T3249;
  wire T3250;
  reg[0:0] dramBank3PortHadValidRequest_1;
  wire T3251;
  wire T3252;
  wire T3253;
  wire T3254;
  wire[4:0] T3255;
  wire T3256;
  wire T3257;
  wire[4:0] T3258;
  wire T3259;
  wire T3260;
  wire T3261;
  wire[9:0] T3262;
  wire T3263;
  wire T3264;
  wire T3265;
  reg[0:0] dramBank2PortHadValidRequest_1;
  wire T3266;
  wire T3267;
  wire T3268;
  wire T3269;
  wire[4:0] T3270;
  wire T3271;
  wire T3272;
  wire[4:0] T3273;
  wire T3274;
  wire T3275;
  wire T3276;
  wire[9:0] T3277;
  wire T3278;
  wire T3279;
  wire T3280;
  reg[0:0] dramBank1PortHadValidRequest_1;
  wire T3281;
  wire T3282;
  wire T3283;
  wire T3284;
  wire[4:0] T3285;
  wire T3286;
  wire T3287;
  wire[4:0] T3288;
  wire T3289;
  wire T3290;
  wire T3291;
  wire[9:0] T3292;
  wire T3293;
  wire T3294;
  reg[0:0] dramBank0PortHadValidRequest_1;
  wire T3295;
  wire T3296;
  wire T3297;
  wire T3298;
  wire[4:0] T3299;
  wire T3300;
  wire T3301;
  wire[4:0] T3302;
  wire T3303;
  wire T3304;
  wire T3305;
  wire[9:0] T3306;
  wire T3307;
  wire T3308;
  wire AllOffloadsValid_0;
  wire T3309;
  wire T3310;
  wire T3311;
  reg[0:0] dramBank7PortHadValidRequest_0;
  wire T3312;
  wire T3313;
  wire T3314;
  wire T3315;
  wire[4:0] T3316;
  wire T3317;
  wire T3318;
  wire[4:0] T3319;
  wire T3320;
  wire T3321;
  wire T3322;
  wire[9:0] T3323;
  wire T3324;
  wire T3325;
  wire T3326;
  reg[0:0] dramBank6PortHadValidRequest_0;
  wire T3327;
  wire T3328;
  wire T3329;
  wire T3330;
  wire[4:0] T3331;
  wire T3332;
  wire T3333;
  wire[4:0] T3334;
  wire T3335;
  wire T3336;
  wire T3337;
  wire[9:0] T3338;
  wire T3339;
  wire T3340;
  wire T3341;
  reg[0:0] dramBank5PortHadValidRequest_0;
  wire T3342;
  wire T3343;
  wire T3344;
  wire T3345;
  wire[4:0] T3346;
  wire T3347;
  wire T3348;
  wire[4:0] T3349;
  wire T3350;
  wire T3351;
  wire T3352;
  wire[9:0] T3353;
  wire T3354;
  wire T3355;
  wire T3356;
  reg[0:0] dramBank4PortHadValidRequest_0;
  wire T3357;
  wire T3358;
  wire T3359;
  wire T3360;
  wire[4:0] T3361;
  wire T3362;
  wire T3363;
  wire[4:0] T3364;
  wire T3365;
  wire T3366;
  wire T3367;
  wire[9:0] T3368;
  wire T3369;
  wire T3370;
  wire T3371;
  reg[0:0] dramBank3PortHadValidRequest_0;
  wire T3372;
  wire T3373;
  wire T3374;
  wire T3375;
  wire[4:0] T3376;
  wire T3377;
  wire T3378;
  wire[4:0] T3379;
  wire T3380;
  wire T3381;
  wire T3382;
  wire[9:0] T3383;
  wire T3384;
  wire T3385;
  wire T3386;
  reg[0:0] dramBank2PortHadValidRequest_0;
  wire T3387;
  wire T3388;
  wire T3389;
  wire T3390;
  wire[4:0] T3391;
  wire T3392;
  wire T3393;
  wire[4:0] T3394;
  wire T3395;
  wire T3396;
  wire T3397;
  wire[9:0] T3398;
  wire T3399;
  wire T3400;
  wire T3401;
  reg[0:0] dramBank1PortHadValidRequest_0;
  wire T3402;
  wire T3403;
  wire T3404;
  wire T3405;
  wire[4:0] T3406;
  wire T3407;
  wire T3408;
  wire[4:0] T3409;
  wire T3410;
  wire T3411;
  wire T3412;
  wire[9:0] T3413;
  wire T3414;
  wire T3415;
  reg[0:0] dramBank0PortHadValidRequest_0;
  wire T3416;
  wire T3417;
  wire T3418;
  wire T3419;
  wire[4:0] T3420;
  wire T3421;
  wire T3422;
  wire[4:0] T3423;
  wire T3424;
  wire T3425;
  wire T3426;
  wire[9:0] T3427;
  wire T3428;
  wire T3429;
  wire T3430;
  wire T3431;
  wire T3432;
  wire T3433;
  wire T3434;
  wire T3435;
  wire T3436;
  wire T3437;
  wire T3438;
  wire T3439;
  wire T3440;
  wire T3441;
  wire T3442;
  wire T3443;
  wire T3444;
  wire T3445;
  wire T3446;
  wire T3447;
  wire T3448;
  wire T3449;
  wire T3450;
  wire T3451;
  wire T3452;
  wire T3453;
  wire T3454;
  wire T3455;
  wire T3456;
  wire T3457;
  wire T3458;
  wire T3459;
  wire T3460;
  wire T3461;
  wire T3462;
  wire T3463;
  wire T3464;
  wire T3465;
  wire[7:0] T3466;
  wire[7:0] T3467;
  wire[7:0] T3468;
  wire[7:0] T3469;
  wire[7:0] T3470;
  wire[7:0] T3471;
  wire[7:0] T3472;
  wire[7:0] T3473;
  wire[7:0] T3474;
  wire[7:0] T3475;
  wire[7:0] T3476;
  wire[7:0] T3477;
  wire[7:0] T3478;
  wire[7:0] T3479;
  wire[7:0] T3480;
  wire[7:0] T3481;
  wire[7:0] T3482;
  wire[7:0] T3483;
  wire[7:0] T3484;
  wire[7:0] T3485;
  wire[7:0] T3486;
  wire[7:0] T3487;
  wire[7:0] T3488;
  wire[7:0] T3489;
  wire[7:0] T3490;
  wire[7:0] T3491;
  wire[7:0] T3492;
  wire[7:0] T3493;
  wire[7:0] T3494;
  wire[7:0] T3495;
  wire[7:0] T3496;
  wire[7:0] T3497;
  wire[7:0] T3498;
  wire[7:0] T3499;
  wire[7:0] T3500;
  wire[7:0] T3501;
  wire[7:0] T3502;
  wire[7:0] T3503;
  wire T3504;
  wire T3505;
  wire T3506;
  wire T3507;
  wire T3508;
  wire T3509;
  wire T3510;
  wire T3511;
  wire T3512;
  wire T3513;
  wire T3514;
  wire T3515;
  wire T3516;
  wire T3517;
  wire T3518;
  wire T3519;
  wire T3520;
  wire T3521;
  wire T3522;
  wire T3523;
  wire T3524;
  wire T3525;
  wire T3526;
  wire T3527;
  wire T3528;
  wire T3529;
  wire T3530;
  wire T3531;
  wire T3532;
  wire T3533;
  wire T3534;
  wire[9:0] T3535;
  wire[9:0] T3536;
  wire[9:0] T3537;
  reg[9:0] inputTag_7;
  wire[9:0] T3538;
  wire[9:0] T3539;
  wire[9:0] T3540;
  wire[9:0] T3541;
  reg[9:0] inputTag_6;
  wire[9:0] T3542;
  wire[9:0] T3543;
  wire[9:0] T3544;
  wire[9:0] T3545;
  reg[9:0] inputTag_5;
  wire[9:0] T3546;
  wire[9:0] T3547;
  wire[9:0] T3548;
  wire[9:0] T3549;
  reg[9:0] inputTag_4;
  wire[9:0] T3550;
  wire[9:0] T3551;
  wire[9:0] T3552;
  wire[9:0] T3553;
  reg[9:0] inputTag_3;
  wire[9:0] T3554;
  wire[9:0] T3555;
  wire[9:0] T3556;
  wire[9:0] T3557;
  reg[9:0] inputTag_2;
  wire[9:0] T3558;
  wire[9:0] T3559;
  wire[9:0] T3560;
  wire[9:0] T3561;
  reg[9:0] inputTag_1;
  wire[9:0] T3562;
  wire[9:0] T3563;
  wire[9:0] T3564;
  reg[9:0] inputTag_0;
  wire[9:0] T3565;
  wire T3566;
  wire T3567;
  wire T3568;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T1 = T3512 && T2;
  assign T2 = State_7 == 8'h0/* 0*/;
  assign T3 = T3430 || T4;
  assign T4 = T765 && T5;
  assign T5 = T6[3'h7/* 7*/];
  assign T6 = T7[3'h7/* 7*/:1'h0/* 0*/];
  assign T7 = 8'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T2581 && AllOffloadsValid_7;
  assign AllOffloadsValid_7 = T9;
  assign T9 = T2477 && T10;
  assign T10 = T2473 || T11;
  assign T11 = ! dramBank7PortHadValidRequest_7;
  assign T12 = T2470 && T13;
  assign T13 = dramBank7PortHadValidRequest_7 || T14;
  assign T14 = T2468 && dramBank7Port_req_valid;
  assign dramBank7Port_req_valid = T15;
  assign T15 = T2385 && T16;
  assign T16 = T2384 && T17;
  assign T17 = T19 == T18;
  assign T18 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T19 = T2364 | T20;
  assign T20 = State_7 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23[3'h7/* 7*/];
  assign T23 = T24[3'h7/* 7*/:1'h0/* 0*/];
  assign T24 = 8'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_7 == 1'h0/* 0*/;
  assign T26 = T30 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_7;
  assign T28 = T29 == vThreadEncoder_io_chosen;
  assign T29 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T30 = T32 && T31;
  assign T31 = State_7 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_7 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = T36 == rThreadEncoder_io_chosen;
  assign T36 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign AllOffloadsReady = T37;
  assign T37 = T49 && T38;
  assign T38 = T45 || T39;
  assign T39 = T41 && T40;
  assign T40 = ! dramBank7Port_req_valid;
  assign T41 = ! dramBank7PortHadReadyRequest;
  assign T42 = T44 && T43;
  assign T43 = dramBank7PortHadReadyRequest || dramBank7Port_req_valid;
  assign T44 = ! AllOffloadsReady;
  assign T45 = dramBank7Port_req_ready || dramBank7_ready_received;
  assign T46 = T48 && T47;
  assign T47 = dramBank7_ready_received || dramBank7Port_req_ready;
  assign dramBank7Port_req_ready = mainOff_dramBank7_req_ready;
  assign mainOff_dramBank7_rep_ready = dramBank7Port_rep_ready;
  assign dramBank7Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank7_req_valid = dramBank7Port_req_valid;
  assign T48 = ! AllOffloadsReady;
  assign T49 = T156 && T50;
  assign T50 = T152 || T51;
  assign T51 = T148 && T52;
  assign T52 = ! dramBank6Port_req_valid;
  assign dramBank6Port_req_valid = T53;
  assign T53 = T58 && T54;
  assign T54 = T57 && T55;
  assign T55 = T19 == T56;
  assign T56 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T57 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T58 = T147 && T59;
  assign T59 = ! T60;
  assign T60 = T71 | T61;
  assign T61 = dramBank6_valid_received_7 & T22;
  assign T62 = T68 && T63;
  assign T63 = dramBank6_valid_received_7 || T64;
  assign T64 = dramBank6Port_rep_valid && T65;
  assign T65 = dramBank6Port_rep_tag == T66;
  assign T66 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank6Port_rep_tag = mainOff_dramBank6_rep_tag;
  assign mainOff_dramBank6_rep_ready = dramBank6Port_rep_ready;
  assign dramBank6Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank6_req_valid = dramBank6Port_req_valid;
  assign mainOff_dramBank6_req_tag = dramBank6Port_req_tag;
  assign dramBank6Port_req_tag = T67;
  assign T67 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank6Port_rep_valid = mainOff_dramBank6_rep_valid;
  assign T68 = ! T69;
  assign T69 = T70 == 5'h7/* 7*/;
  assign T70 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T71 = T82 | T72;
  assign T72 = dramBank6_valid_received_6 & T73;
  assign T73 = T23[3'h6/* 6*/];
  assign T74 = T79 && T75;
  assign T75 = dramBank6_valid_received_6 || T76;
  assign T76 = dramBank6Port_rep_valid && T77;
  assign T77 = dramBank6Port_rep_tag == T78;
  assign T78 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T79 = ! T80;
  assign T80 = T81 == 5'h6/* 6*/;
  assign T81 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T82 = T93 | T83;
  assign T83 = dramBank6_valid_received_5 & T84;
  assign T84 = T23[3'h5/* 5*/];
  assign T85 = T90 && T86;
  assign T86 = dramBank6_valid_received_5 || T87;
  assign T87 = dramBank6Port_rep_valid && T88;
  assign T88 = dramBank6Port_rep_tag == T89;
  assign T89 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T90 = ! T91;
  assign T91 = T92 == 5'h5/* 5*/;
  assign T92 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T93 = T104 | T94;
  assign T94 = dramBank6_valid_received_4 & T95;
  assign T95 = T23[3'h4/* 4*/];
  assign T96 = T101 && T97;
  assign T97 = dramBank6_valid_received_4 || T98;
  assign T98 = dramBank6Port_rep_valid && T99;
  assign T99 = dramBank6Port_rep_tag == T100;
  assign T100 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T101 = ! T102;
  assign T102 = T103 == 5'h4/* 4*/;
  assign T103 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T104 = T115 | T105;
  assign T105 = dramBank6_valid_received_3 & T106;
  assign T106 = T23[2'h3/* 3*/];
  assign T107 = T112 && T108;
  assign T108 = dramBank6_valid_received_3 || T109;
  assign T109 = dramBank6Port_rep_valid && T110;
  assign T110 = dramBank6Port_rep_tag == T111;
  assign T111 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T112 = ! T113;
  assign T113 = T114 == 5'h3/* 3*/;
  assign T114 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T115 = T126 | T116;
  assign T116 = dramBank6_valid_received_2 & T117;
  assign T117 = T23[2'h2/* 2*/];
  assign T118 = T123 && T119;
  assign T119 = dramBank6_valid_received_2 || T120;
  assign T120 = dramBank6Port_rep_valid && T121;
  assign T121 = dramBank6Port_rep_tag == T122;
  assign T122 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T123 = ! T124;
  assign T124 = T125 == 5'h2/* 2*/;
  assign T125 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T126 = T137 | T127;
  assign T127 = dramBank6_valid_received_1 & T128;
  assign T128 = T23[1'h1/* 1*/];
  assign T129 = T134 && T130;
  assign T130 = dramBank6_valid_received_1 || T131;
  assign T131 = dramBank6Port_rep_valid && T132;
  assign T132 = dramBank6Port_rep_tag == T133;
  assign T133 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T134 = ! T135;
  assign T135 = T136 == 5'h1/* 1*/;
  assign T136 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T137 = dramBank6_valid_received_0 & T138;
  assign T138 = T23[1'h0/* 0*/];
  assign T139 = T144 && T140;
  assign T140 = dramBank6_valid_received_0 || T141;
  assign T141 = dramBank6Port_rep_valid && T142;
  assign T142 = dramBank6Port_rep_tag == T143;
  assign T143 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T148 = ! dramBank6PortHadReadyRequest;
  assign T149 = T151 && T150;
  assign T150 = dramBank6PortHadReadyRequest || dramBank6Port_req_valid;
  assign T151 = ! AllOffloadsReady;
  assign T152 = dramBank6Port_req_ready || dramBank6_ready_received;
  assign T153 = T155 && T154;
  assign T154 = dramBank6_ready_received || dramBank6Port_req_ready;
  assign dramBank6Port_req_ready = mainOff_dramBank6_req_ready;
  assign T155 = ! AllOffloadsReady;
  assign T156 = T256 && T157;
  assign T157 = T252 || T158;
  assign T158 = T248 && T159;
  assign T159 = ! dramBank5Port_req_valid;
  assign dramBank5Port_req_valid = T160;
  assign T160 = T165 && T161;
  assign T161 = T164 && T162;
  assign T162 = T19 == T163;
  assign T163 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T164 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T165 = T247 && T166;
  assign T166 = ! T167;
  assign T167 = T178 | T168;
  assign T168 = dramBank5_valid_received_7 & T22;
  assign T169 = T175 && T170;
  assign T170 = dramBank5_valid_received_7 || T171;
  assign T171 = dramBank5Port_rep_valid && T172;
  assign T172 = dramBank5Port_rep_tag == T173;
  assign T173 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank5Port_rep_tag = mainOff_dramBank5_rep_tag;
  assign mainOff_dramBank5_rep_ready = dramBank5Port_rep_ready;
  assign dramBank5Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank5_req_valid = dramBank5Port_req_valid;
  assign mainOff_dramBank5_req_tag = dramBank5Port_req_tag;
  assign dramBank5Port_req_tag = T174;
  assign T174 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank5Port_rep_valid = mainOff_dramBank5_rep_valid;
  assign T175 = ! T176;
  assign T176 = T177 == 5'h7/* 7*/;
  assign T177 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T178 = T188 | T179;
  assign T179 = dramBank5_valid_received_6 & T73;
  assign T180 = T185 && T181;
  assign T181 = dramBank5_valid_received_6 || T182;
  assign T182 = dramBank5Port_rep_valid && T183;
  assign T183 = dramBank5Port_rep_tag == T184;
  assign T184 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T185 = ! T186;
  assign T186 = T187 == 5'h6/* 6*/;
  assign T187 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T188 = T198 | T189;
  assign T189 = dramBank5_valid_received_5 & T84;
  assign T190 = T195 && T191;
  assign T191 = dramBank5_valid_received_5 || T192;
  assign T192 = dramBank5Port_rep_valid && T193;
  assign T193 = dramBank5Port_rep_tag == T194;
  assign T194 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T195 = ! T196;
  assign T196 = T197 == 5'h5/* 5*/;
  assign T197 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T198 = T208 | T199;
  assign T199 = dramBank5_valid_received_4 & T95;
  assign T200 = T205 && T201;
  assign T201 = dramBank5_valid_received_4 || T202;
  assign T202 = dramBank5Port_rep_valid && T203;
  assign T203 = dramBank5Port_rep_tag == T204;
  assign T204 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T205 = ! T206;
  assign T206 = T207 == 5'h4/* 4*/;
  assign T207 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T208 = T218 | T209;
  assign T209 = dramBank5_valid_received_3 & T106;
  assign T210 = T215 && T211;
  assign T211 = dramBank5_valid_received_3 || T212;
  assign T212 = dramBank5Port_rep_valid && T213;
  assign T213 = dramBank5Port_rep_tag == T214;
  assign T214 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T215 = ! T216;
  assign T216 = T217 == 5'h3/* 3*/;
  assign T217 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T218 = T228 | T219;
  assign T219 = dramBank5_valid_received_2 & T117;
  assign T220 = T225 && T221;
  assign T221 = dramBank5_valid_received_2 || T222;
  assign T222 = dramBank5Port_rep_valid && T223;
  assign T223 = dramBank5Port_rep_tag == T224;
  assign T224 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T225 = ! T226;
  assign T226 = T227 == 5'h2/* 2*/;
  assign T227 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T228 = T238 | T229;
  assign T229 = dramBank5_valid_received_1 & T128;
  assign T230 = T235 && T231;
  assign T231 = dramBank5_valid_received_1 || T232;
  assign T232 = dramBank5Port_rep_valid && T233;
  assign T233 = dramBank5Port_rep_tag == T234;
  assign T234 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T235 = ! T236;
  assign T236 = T237 == 5'h1/* 1*/;
  assign T237 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T238 = dramBank5_valid_received_0 & T138;
  assign T239 = T244 && T240;
  assign T240 = dramBank5_valid_received_0 || T241;
  assign T241 = dramBank5Port_rep_valid && T242;
  assign T242 = dramBank5Port_rep_tag == T243;
  assign T243 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T244 = ! T245;
  assign T245 = T246 == 5'h0/* 0*/;
  assign T246 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T247 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T248 = ! dramBank5PortHadReadyRequest;
  assign T249 = T251 && T250;
  assign T250 = dramBank5PortHadReadyRequest || dramBank5Port_req_valid;
  assign T251 = ! AllOffloadsReady;
  assign T252 = dramBank5Port_req_ready || dramBank5_ready_received;
  assign T253 = T255 && T254;
  assign T254 = dramBank5_ready_received || dramBank5Port_req_ready;
  assign dramBank5Port_req_ready = mainOff_dramBank5_req_ready;
  assign T255 = ! AllOffloadsReady;
  assign T256 = T356 && T257;
  assign T257 = T352 || T258;
  assign T258 = T348 && T259;
  assign T259 = ! dramBank4Port_req_valid;
  assign dramBank4Port_req_valid = T260;
  assign T260 = T265 && T261;
  assign T261 = T264 && T262;
  assign T262 = T19 == T263;
  assign T263 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T264 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T265 = T347 && T266;
  assign T266 = ! T267;
  assign T267 = T278 | T268;
  assign T268 = dramBank4_valid_received_7 & T22;
  assign T269 = T275 && T270;
  assign T270 = dramBank4_valid_received_7 || T271;
  assign T271 = dramBank4Port_rep_valid && T272;
  assign T272 = dramBank4Port_rep_tag == T273;
  assign T273 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank4Port_rep_tag = mainOff_dramBank4_rep_tag;
  assign mainOff_dramBank4_rep_ready = dramBank4Port_rep_ready;
  assign dramBank4Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank4_req_valid = dramBank4Port_req_valid;
  assign mainOff_dramBank4_req_tag = dramBank4Port_req_tag;
  assign dramBank4Port_req_tag = T274;
  assign T274 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank4Port_rep_valid = mainOff_dramBank4_rep_valid;
  assign T275 = ! T276;
  assign T276 = T277 == 5'h7/* 7*/;
  assign T277 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T278 = T288 | T279;
  assign T279 = dramBank4_valid_received_6 & T73;
  assign T280 = T285 && T281;
  assign T281 = dramBank4_valid_received_6 || T282;
  assign T282 = dramBank4Port_rep_valid && T283;
  assign T283 = dramBank4Port_rep_tag == T284;
  assign T284 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T285 = ! T286;
  assign T286 = T287 == 5'h6/* 6*/;
  assign T287 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T288 = T298 | T289;
  assign T289 = dramBank4_valid_received_5 & T84;
  assign T290 = T295 && T291;
  assign T291 = dramBank4_valid_received_5 || T292;
  assign T292 = dramBank4Port_rep_valid && T293;
  assign T293 = dramBank4Port_rep_tag == T294;
  assign T294 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T295 = ! T296;
  assign T296 = T297 == 5'h5/* 5*/;
  assign T297 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T298 = T308 | T299;
  assign T299 = dramBank4_valid_received_4 & T95;
  assign T300 = T305 && T301;
  assign T301 = dramBank4_valid_received_4 || T302;
  assign T302 = dramBank4Port_rep_valid && T303;
  assign T303 = dramBank4Port_rep_tag == T304;
  assign T304 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T305 = ! T306;
  assign T306 = T307 == 5'h4/* 4*/;
  assign T307 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T308 = T318 | T309;
  assign T309 = dramBank4_valid_received_3 & T106;
  assign T310 = T315 && T311;
  assign T311 = dramBank4_valid_received_3 || T312;
  assign T312 = dramBank4Port_rep_valid && T313;
  assign T313 = dramBank4Port_rep_tag == T314;
  assign T314 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T315 = ! T316;
  assign T316 = T317 == 5'h3/* 3*/;
  assign T317 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T318 = T328 | T319;
  assign T319 = dramBank4_valid_received_2 & T117;
  assign T320 = T325 && T321;
  assign T321 = dramBank4_valid_received_2 || T322;
  assign T322 = dramBank4Port_rep_valid && T323;
  assign T323 = dramBank4Port_rep_tag == T324;
  assign T324 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T325 = ! T326;
  assign T326 = T327 == 5'h2/* 2*/;
  assign T327 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T328 = T338 | T329;
  assign T329 = dramBank4_valid_received_1 & T128;
  assign T330 = T335 && T331;
  assign T331 = dramBank4_valid_received_1 || T332;
  assign T332 = dramBank4Port_rep_valid && T333;
  assign T333 = dramBank4Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T335 = ! T336;
  assign T336 = T337 == 5'h1/* 1*/;
  assign T337 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T338 = dramBank4_valid_received_0 & T138;
  assign T339 = T344 && T340;
  assign T340 = dramBank4_valid_received_0 || T341;
  assign T341 = dramBank4Port_rep_valid && T342;
  assign T342 = dramBank4Port_rep_tag == T343;
  assign T343 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T344 = ! T345;
  assign T345 = T346 == 5'h0/* 0*/;
  assign T346 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T347 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T348 = ! dramBank4PortHadReadyRequest;
  assign T349 = T351 && T350;
  assign T350 = dramBank4PortHadReadyRequest || dramBank4Port_req_valid;
  assign T351 = ! AllOffloadsReady;
  assign T352 = dramBank4Port_req_ready || dramBank4_ready_received;
  assign T353 = T355 && T354;
  assign T354 = dramBank4_ready_received || dramBank4Port_req_ready;
  assign dramBank4Port_req_ready = mainOff_dramBank4_req_ready;
  assign T355 = ! AllOffloadsReady;
  assign T356 = T456 && T357;
  assign T357 = T452 || T358;
  assign T358 = T448 && T359;
  assign T359 = ! dramBank3Port_req_valid;
  assign dramBank3Port_req_valid = T360;
  assign T360 = T365 && T361;
  assign T361 = T364 && T362;
  assign T362 = T19 == T363;
  assign T363 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T364 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T365 = T447 && T366;
  assign T366 = ! T367;
  assign T367 = T378 | T368;
  assign T368 = dramBank3_valid_received_7 & T22;
  assign T369 = T375 && T370;
  assign T370 = dramBank3_valid_received_7 || T371;
  assign T371 = dramBank3Port_rep_valid && T372;
  assign T372 = dramBank3Port_rep_tag == T373;
  assign T373 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank3Port_rep_tag = mainOff_dramBank3_rep_tag;
  assign mainOff_dramBank3_rep_ready = dramBank3Port_rep_ready;
  assign dramBank3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank3_req_valid = dramBank3Port_req_valid;
  assign mainOff_dramBank3_req_tag = dramBank3Port_req_tag;
  assign dramBank3Port_req_tag = T374;
  assign T374 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank3Port_rep_valid = mainOff_dramBank3_rep_valid;
  assign T375 = ! T376;
  assign T376 = T377 == 5'h7/* 7*/;
  assign T377 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T378 = T388 | T379;
  assign T379 = dramBank3_valid_received_6 & T73;
  assign T380 = T385 && T381;
  assign T381 = dramBank3_valid_received_6 || T382;
  assign T382 = dramBank3Port_rep_valid && T383;
  assign T383 = dramBank3Port_rep_tag == T384;
  assign T384 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T385 = ! T386;
  assign T386 = T387 == 5'h6/* 6*/;
  assign T387 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T388 = T398 | T389;
  assign T389 = dramBank3_valid_received_5 & T84;
  assign T390 = T395 && T391;
  assign T391 = dramBank3_valid_received_5 || T392;
  assign T392 = dramBank3Port_rep_valid && T393;
  assign T393 = dramBank3Port_rep_tag == T394;
  assign T394 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T395 = ! T396;
  assign T396 = T397 == 5'h5/* 5*/;
  assign T397 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T398 = T408 | T399;
  assign T399 = dramBank3_valid_received_4 & T95;
  assign T400 = T405 && T401;
  assign T401 = dramBank3_valid_received_4 || T402;
  assign T402 = dramBank3Port_rep_valid && T403;
  assign T403 = dramBank3Port_rep_tag == T404;
  assign T404 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T405 = ! T406;
  assign T406 = T407 == 5'h4/* 4*/;
  assign T407 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T408 = T418 | T409;
  assign T409 = dramBank3_valid_received_3 & T106;
  assign T410 = T415 && T411;
  assign T411 = dramBank3_valid_received_3 || T412;
  assign T412 = dramBank3Port_rep_valid && T413;
  assign T413 = dramBank3Port_rep_tag == T414;
  assign T414 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T415 = ! T416;
  assign T416 = T417 == 5'h3/* 3*/;
  assign T417 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T418 = T428 | T419;
  assign T419 = dramBank3_valid_received_2 & T117;
  assign T420 = T425 && T421;
  assign T421 = dramBank3_valid_received_2 || T422;
  assign T422 = dramBank3Port_rep_valid && T423;
  assign T423 = dramBank3Port_rep_tag == T424;
  assign T424 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T425 = ! T426;
  assign T426 = T427 == 5'h2/* 2*/;
  assign T427 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T428 = T438 | T429;
  assign T429 = dramBank3_valid_received_1 & T128;
  assign T430 = T435 && T431;
  assign T431 = dramBank3_valid_received_1 || T432;
  assign T432 = dramBank3Port_rep_valid && T433;
  assign T433 = dramBank3Port_rep_tag == T434;
  assign T434 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T435 = ! T436;
  assign T436 = T437 == 5'h1/* 1*/;
  assign T437 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T438 = dramBank3_valid_received_0 & T138;
  assign T439 = T444 && T440;
  assign T440 = dramBank3_valid_received_0 || T441;
  assign T441 = dramBank3Port_rep_valid && T442;
  assign T442 = dramBank3Port_rep_tag == T443;
  assign T443 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T444 = ! T445;
  assign T445 = T446 == 5'h0/* 0*/;
  assign T446 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T447 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T448 = ! dramBank3PortHadReadyRequest;
  assign T449 = T451 && T450;
  assign T450 = dramBank3PortHadReadyRequest || dramBank3Port_req_valid;
  assign T451 = ! AllOffloadsReady;
  assign T452 = dramBank3Port_req_ready || dramBank3_ready_received;
  assign T453 = T455 && T454;
  assign T454 = dramBank3_ready_received || dramBank3Port_req_ready;
  assign dramBank3Port_req_ready = mainOff_dramBank3_req_ready;
  assign T455 = ! AllOffloadsReady;
  assign T456 = T556 && T457;
  assign T457 = T552 || T458;
  assign T458 = T548 && T459;
  assign T459 = ! dramBank2Port_req_valid;
  assign dramBank2Port_req_valid = T460;
  assign T460 = T465 && T461;
  assign T461 = T464 && T462;
  assign T462 = T19 == T463;
  assign T463 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T464 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T465 = T547 && T466;
  assign T466 = ! T467;
  assign T467 = T478 | T468;
  assign T468 = dramBank2_valid_received_7 & T22;
  assign T469 = T475 && T470;
  assign T470 = dramBank2_valid_received_7 || T471;
  assign T471 = dramBank2Port_rep_valid && T472;
  assign T472 = dramBank2Port_rep_tag == T473;
  assign T473 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank2Port_rep_tag = mainOff_dramBank2_rep_tag;
  assign mainOff_dramBank2_rep_ready = dramBank2Port_rep_ready;
  assign dramBank2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank2_req_valid = dramBank2Port_req_valid;
  assign mainOff_dramBank2_req_tag = dramBank2Port_req_tag;
  assign dramBank2Port_req_tag = T474;
  assign T474 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank2Port_rep_valid = mainOff_dramBank2_rep_valid;
  assign T475 = ! T476;
  assign T476 = T477 == 5'h7/* 7*/;
  assign T477 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T478 = T488 | T479;
  assign T479 = dramBank2_valid_received_6 & T73;
  assign T480 = T485 && T481;
  assign T481 = dramBank2_valid_received_6 || T482;
  assign T482 = dramBank2Port_rep_valid && T483;
  assign T483 = dramBank2Port_rep_tag == T484;
  assign T484 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T485 = ! T486;
  assign T486 = T487 == 5'h6/* 6*/;
  assign T487 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T488 = T498 | T489;
  assign T489 = dramBank2_valid_received_5 & T84;
  assign T490 = T495 && T491;
  assign T491 = dramBank2_valid_received_5 || T492;
  assign T492 = dramBank2Port_rep_valid && T493;
  assign T493 = dramBank2Port_rep_tag == T494;
  assign T494 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T495 = ! T496;
  assign T496 = T497 == 5'h5/* 5*/;
  assign T497 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T498 = T508 | T499;
  assign T499 = dramBank2_valid_received_4 & T95;
  assign T500 = T505 && T501;
  assign T501 = dramBank2_valid_received_4 || T502;
  assign T502 = dramBank2Port_rep_valid && T503;
  assign T503 = dramBank2Port_rep_tag == T504;
  assign T504 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T505 = ! T506;
  assign T506 = T507 == 5'h4/* 4*/;
  assign T507 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T508 = T518 | T509;
  assign T509 = dramBank2_valid_received_3 & T106;
  assign T510 = T515 && T511;
  assign T511 = dramBank2_valid_received_3 || T512;
  assign T512 = dramBank2Port_rep_valid && T513;
  assign T513 = dramBank2Port_rep_tag == T514;
  assign T514 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T515 = ! T516;
  assign T516 = T517 == 5'h3/* 3*/;
  assign T517 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T518 = T528 | T519;
  assign T519 = dramBank2_valid_received_2 & T117;
  assign T520 = T525 && T521;
  assign T521 = dramBank2_valid_received_2 || T522;
  assign T522 = dramBank2Port_rep_valid && T523;
  assign T523 = dramBank2Port_rep_tag == T524;
  assign T524 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T525 = ! T526;
  assign T526 = T527 == 5'h2/* 2*/;
  assign T527 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T528 = T538 | T529;
  assign T529 = dramBank2_valid_received_1 & T128;
  assign T530 = T535 && T531;
  assign T531 = dramBank2_valid_received_1 || T532;
  assign T532 = dramBank2Port_rep_valid && T533;
  assign T533 = dramBank2Port_rep_tag == T534;
  assign T534 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T535 = ! T536;
  assign T536 = T537 == 5'h1/* 1*/;
  assign T537 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T538 = dramBank2_valid_received_0 & T138;
  assign T539 = T544 && T540;
  assign T540 = dramBank2_valid_received_0 || T541;
  assign T541 = dramBank2Port_rep_valid && T542;
  assign T542 = dramBank2Port_rep_tag == T543;
  assign T543 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T544 = ! T545;
  assign T545 = T546 == 5'h0/* 0*/;
  assign T546 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T547 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T548 = ! dramBank2PortHadReadyRequest;
  assign T549 = T551 && T550;
  assign T550 = dramBank2PortHadReadyRequest || dramBank2Port_req_valid;
  assign T551 = ! AllOffloadsReady;
  assign T552 = dramBank2Port_req_ready || dramBank2_ready_received;
  assign T553 = T555 && T554;
  assign T554 = dramBank2_ready_received || dramBank2Port_req_ready;
  assign dramBank2Port_req_ready = mainOff_dramBank2_req_ready;
  assign T555 = ! AllOffloadsReady;
  assign T556 = T656 && T557;
  assign T557 = T652 || T558;
  assign T558 = T648 && T559;
  assign T559 = ! dramBank1Port_req_valid;
  assign dramBank1Port_req_valid = T560;
  assign T560 = T565 && T561;
  assign T561 = T564 && T562;
  assign T562 = T19 == T563;
  assign T563 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T564 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T565 = T647 && T566;
  assign T566 = ! T567;
  assign T567 = T578 | T568;
  assign T568 = dramBank1_valid_received_7 & T22;
  assign T569 = T575 && T570;
  assign T570 = dramBank1_valid_received_7 || T571;
  assign T571 = dramBank1Port_rep_valid && T572;
  assign T572 = dramBank1Port_rep_tag == T573;
  assign T573 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank1Port_rep_tag = mainOff_dramBank1_rep_tag;
  assign mainOff_dramBank1_rep_ready = dramBank1Port_rep_ready;
  assign dramBank1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank1_req_valid = dramBank1Port_req_valid;
  assign mainOff_dramBank1_req_tag = dramBank1Port_req_tag;
  assign dramBank1Port_req_tag = T574;
  assign T574 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank1Port_rep_valid = mainOff_dramBank1_rep_valid;
  assign T575 = ! T576;
  assign T576 = T577 == 5'h7/* 7*/;
  assign T577 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T578 = T588 | T579;
  assign T579 = dramBank1_valid_received_6 & T73;
  assign T580 = T585 && T581;
  assign T581 = dramBank1_valid_received_6 || T582;
  assign T582 = dramBank1Port_rep_valid && T583;
  assign T583 = dramBank1Port_rep_tag == T584;
  assign T584 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T585 = ! T586;
  assign T586 = T587 == 5'h6/* 6*/;
  assign T587 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T588 = T598 | T589;
  assign T589 = dramBank1_valid_received_5 & T84;
  assign T590 = T595 && T591;
  assign T591 = dramBank1_valid_received_5 || T592;
  assign T592 = dramBank1Port_rep_valid && T593;
  assign T593 = dramBank1Port_rep_tag == T594;
  assign T594 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T595 = ! T596;
  assign T596 = T597 == 5'h5/* 5*/;
  assign T597 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T598 = T608 | T599;
  assign T599 = dramBank1_valid_received_4 & T95;
  assign T600 = T605 && T601;
  assign T601 = dramBank1_valid_received_4 || T602;
  assign T602 = dramBank1Port_rep_valid && T603;
  assign T603 = dramBank1Port_rep_tag == T604;
  assign T604 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T605 = ! T606;
  assign T606 = T607 == 5'h4/* 4*/;
  assign T607 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T608 = T618 | T609;
  assign T609 = dramBank1_valid_received_3 & T106;
  assign T610 = T615 && T611;
  assign T611 = dramBank1_valid_received_3 || T612;
  assign T612 = dramBank1Port_rep_valid && T613;
  assign T613 = dramBank1Port_rep_tag == T614;
  assign T614 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T615 = ! T616;
  assign T616 = T617 == 5'h3/* 3*/;
  assign T617 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T618 = T628 | T619;
  assign T619 = dramBank1_valid_received_2 & T117;
  assign T620 = T625 && T621;
  assign T621 = dramBank1_valid_received_2 || T622;
  assign T622 = dramBank1Port_rep_valid && T623;
  assign T623 = dramBank1Port_rep_tag == T624;
  assign T624 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T625 = ! T626;
  assign T626 = T627 == 5'h2/* 2*/;
  assign T627 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T628 = T638 | T629;
  assign T629 = dramBank1_valid_received_1 & T128;
  assign T630 = T635 && T631;
  assign T631 = dramBank1_valid_received_1 || T632;
  assign T632 = dramBank1Port_rep_valid && T633;
  assign T633 = dramBank1Port_rep_tag == T634;
  assign T634 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T635 = ! T636;
  assign T636 = T637 == 5'h1/* 1*/;
  assign T637 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T638 = dramBank1_valid_received_0 & T138;
  assign T639 = T644 && T640;
  assign T640 = dramBank1_valid_received_0 || T641;
  assign T641 = dramBank1Port_rep_valid && T642;
  assign T642 = dramBank1Port_rep_tag == T643;
  assign T643 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T644 = ! T645;
  assign T645 = T646 == 5'h0/* 0*/;
  assign T646 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T647 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T648 = ! dramBank1PortHadReadyRequest;
  assign T649 = T651 && T650;
  assign T650 = dramBank1PortHadReadyRequest || dramBank1Port_req_valid;
  assign T651 = ! AllOffloadsReady;
  assign T652 = dramBank1Port_req_ready || dramBank1_ready_received;
  assign T653 = T655 && T654;
  assign T654 = dramBank1_ready_received || dramBank1Port_req_ready;
  assign dramBank1Port_req_ready = mainOff_dramBank1_req_ready;
  assign T655 = ! AllOffloadsReady;
  assign T656 = T751 || T657;
  assign T657 = T747 && T658;
  assign T658 = ! dramBank0Port_req_valid;
  assign dramBank0Port_req_valid = T659;
  assign T659 = T664 && T660;
  assign T660 = T663 && T661;
  assign T661 = T19 == T662;
  assign T662 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T663 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T664 = T746 && T665;
  assign T665 = ! T666;
  assign T666 = T677 | T667;
  assign T667 = dramBank0_valid_received_7 & T22;
  assign T668 = T674 && T669;
  assign T669 = dramBank0_valid_received_7 || T670;
  assign T670 = dramBank0Port_rep_valid && T671;
  assign T671 = dramBank0Port_rep_tag == T672;
  assign T672 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank0Port_rep_tag = mainOff_dramBank0_rep_tag;
  assign mainOff_dramBank0_rep_ready = dramBank0Port_rep_ready;
  assign dramBank0Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank0_req_valid = dramBank0Port_req_valid;
  assign mainOff_dramBank0_req_tag = dramBank0Port_req_tag;
  assign dramBank0Port_req_tag = T673;
  assign T673 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank0Port_rep_valid = mainOff_dramBank0_rep_valid;
  assign T674 = ! T675;
  assign T675 = T676 == 5'h7/* 7*/;
  assign T676 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T677 = T687 | T678;
  assign T678 = dramBank0_valid_received_6 & T73;
  assign T679 = T684 && T680;
  assign T680 = dramBank0_valid_received_6 || T681;
  assign T681 = dramBank0Port_rep_valid && T682;
  assign T682 = dramBank0Port_rep_tag == T683;
  assign T683 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T684 = ! T685;
  assign T685 = T686 == 5'h6/* 6*/;
  assign T686 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T687 = T697 | T688;
  assign T688 = dramBank0_valid_received_5 & T84;
  assign T689 = T694 && T690;
  assign T690 = dramBank0_valid_received_5 || T691;
  assign T691 = dramBank0Port_rep_valid && T692;
  assign T692 = dramBank0Port_rep_tag == T693;
  assign T693 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T694 = ! T695;
  assign T695 = T696 == 5'h5/* 5*/;
  assign T696 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T697 = T707 | T698;
  assign T698 = dramBank0_valid_received_4 & T95;
  assign T699 = T704 && T700;
  assign T700 = dramBank0_valid_received_4 || T701;
  assign T701 = dramBank0Port_rep_valid && T702;
  assign T702 = dramBank0Port_rep_tag == T703;
  assign T703 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T704 = ! T705;
  assign T705 = T706 == 5'h4/* 4*/;
  assign T706 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T707 = T717 | T708;
  assign T708 = dramBank0_valid_received_3 & T106;
  assign T709 = T714 && T710;
  assign T710 = dramBank0_valid_received_3 || T711;
  assign T711 = dramBank0Port_rep_valid && T712;
  assign T712 = dramBank0Port_rep_tag == T713;
  assign T713 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h3/* 3*/;
  assign T716 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T727 | T718;
  assign T718 = dramBank0_valid_received_2 & T117;
  assign T719 = T724 && T720;
  assign T720 = dramBank0_valid_received_2 || T721;
  assign T721 = dramBank0Port_rep_valid && T722;
  assign T722 = dramBank0Port_rep_tag == T723;
  assign T723 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T724 = ! T725;
  assign T725 = T726 == 5'h2/* 2*/;
  assign T726 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T727 = T737 | T728;
  assign T728 = dramBank0_valid_received_1 & T128;
  assign T729 = T734 && T730;
  assign T730 = dramBank0_valid_received_1 || T731;
  assign T731 = dramBank0Port_rep_valid && T732;
  assign T732 = dramBank0Port_rep_tag == T733;
  assign T733 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T734 = ! T735;
  assign T735 = T736 == 5'h1/* 1*/;
  assign T736 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T737 = dramBank0_valid_received_0 & T138;
  assign T738 = T743 && T739;
  assign T739 = dramBank0_valid_received_0 || T740;
  assign T740 = dramBank0Port_rep_valid && T741;
  assign T741 = dramBank0Port_rep_tag == T742;
  assign T742 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h0/* 0*/;
  assign T745 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T747 = ! dramBank0PortHadReadyRequest;
  assign T748 = T750 && T749;
  assign T749 = dramBank0PortHadReadyRequest || dramBank0Port_req_valid;
  assign T750 = ! AllOffloadsReady;
  assign T751 = dramBank0Port_req_ready || dramBank0_ready_received;
  assign T752 = T754 && T753;
  assign T753 = dramBank0_ready_received || dramBank0Port_req_ready;
  assign dramBank0Port_req_ready = mainOff_dramBank0_req_ready;
  assign T754 = ! AllOffloadsReady;
  assign T755 = subStateTh_6 == 1'h0/* 0*/;
  assign T756 = T760 ? 1'h1/* 1*/ : T757;
  assign T757 = T758 ? 1'h0/* 0*/ : subStateTh_6;
  assign T758 = T759 == vThreadEncoder_io_chosen;
  assign T759 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T760 = T2286 && T761;
  assign T761 = State_6 != 8'hff/* 255*/;
  assign T762 = T2204 || T763;
  assign T763 = T765 && T764;
  assign T764 = T6[3'h6/* 6*/];
  assign T765 = T2203 && T766;
  assign T766 = T768 == T767;
  assign T767 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T768 = T771 | T769;
  assign T769 = State_7 & T770;
  assign T770 = {4'h8/* 8*/{T5}};
  assign T771 = T774 | T772;
  assign T772 = State_6 & T773;
  assign T773 = {4'h8/* 8*/{T764}};
  assign T774 = T1774 | T775;
  assign T775 = State_5 & T776;
  assign T776 = {4'h8/* 8*/{T777}};
  assign T777 = T6[3'h5/* 5*/];
  assign T778 = T780 || T779;
  assign T779 = T765 && T777;
  assign T780 = T786 || T781;
  assign T781 = T782 && T777;
  assign T782 = T785 && T783;
  assign T783 = T768 == T784;
  assign T784 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T785 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T786 = T792 || T787;
  assign T787 = T788 && T777;
  assign T788 = T791 && T789;
  assign T789 = T768 == T790;
  assign T790 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T791 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T792 = T798 || T793;
  assign T793 = T794 && T777;
  assign T794 = T797 && T795;
  assign T795 = T768 == T796;
  assign T796 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T797 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T798 = T804 || T799;
  assign T799 = T800 && T777;
  assign T800 = T803 && T801;
  assign T801 = T768 == T802;
  assign T802 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T803 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T804 = T810 || T805;
  assign T805 = T806 && T777;
  assign T806 = T809 && T807;
  assign T807 = T768 == T808;
  assign T808 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T809 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T810 = T816 || T811;
  assign T811 = T812 && T777;
  assign T812 = T815 && T813;
  assign T813 = T768 == T814;
  assign T814 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T815 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T816 = T822 || T817;
  assign T817 = T818 && T777;
  assign T818 = T821 && T819;
  assign T819 = T768 == T820;
  assign T820 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T821 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T822 = T828 || T823;
  assign T823 = T824 && T777;
  assign T824 = T827 && T825;
  assign T825 = T768 == T826;
  assign T826 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T827 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T828 = T924 || T829;
  assign T829 = T830 && T777;
  assign T830 = T892 && T831;
  assign T831 = ! T832;
  assign T832 = b == T833;
  assign T833 = {16'h0/* 0*/, 32'h7/* 7*/};
  assign b = T834 & 48'h7fff/* 32767*/;
  assign T834 = {16'h0/* 0*/, T835};
  assign T835 = T836 >> 33'hc/* 12*/;
  assign T836 = T846 | T837;
  assign T837 = inputReg_7_addr & T838;
  assign T838 = {6'h20/* 32*/{T5}};
  assign T839 = T843 && T840;
  assign T840 = T841[3'h7/* 7*/];
  assign T841 = T842[3'h7/* 7*/:1'h0/* 0*/];
  assign T842 = 8'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T843 = T844 && io_in_valid;
  assign T844 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T845 = T839 ? io_in_bits_addr : inputReg_7_addr;
  assign T846 = T852 | T847;
  assign T847 = inputReg_6_addr & T848;
  assign T848 = {6'h20/* 32*/{T764}};
  assign T849 = T843 && T850;
  assign T850 = T841[3'h6/* 6*/];
  assign T851 = T849 ? io_in_bits_addr : inputReg_6_addr;
  assign T852 = T858 | T853;
  assign T853 = inputReg_5_addr & T854;
  assign T854 = {6'h20/* 32*/{T777}};
  assign T855 = T843 && T856;
  assign T856 = T841[3'h5/* 5*/];
  assign T857 = T855 ? io_in_bits_addr : inputReg_5_addr;
  assign T858 = T865 | T859;
  assign T859 = inputReg_4_addr & T860;
  assign T860 = {6'h20/* 32*/{T861}};
  assign T861 = T6[3'h4/* 4*/];
  assign T862 = T843 && T863;
  assign T863 = T841[3'h4/* 4*/];
  assign T864 = T862 ? io_in_bits_addr : inputReg_4_addr;
  assign T865 = T872 | T866;
  assign T866 = inputReg_3_addr & T867;
  assign T867 = {6'h20/* 32*/{T868}};
  assign T868 = T6[2'h3/* 3*/];
  assign T869 = T843 && T870;
  assign T870 = T841[2'h3/* 3*/];
  assign T871 = T869 ? io_in_bits_addr : inputReg_3_addr;
  assign T872 = T879 | T873;
  assign T873 = inputReg_2_addr & T874;
  assign T874 = {6'h20/* 32*/{T875}};
  assign T875 = T6[2'h2/* 2*/];
  assign T876 = T843 && T877;
  assign T877 = T841[2'h2/* 2*/];
  assign T878 = T876 ? io_in_bits_addr : inputReg_2_addr;
  assign T879 = T886 | T880;
  assign T880 = inputReg_1_addr & T881;
  assign T881 = {6'h20/* 32*/{T882}};
  assign T882 = T6[1'h1/* 1*/];
  assign T883 = T843 && T884;
  assign T884 = T841[1'h1/* 1*/];
  assign T885 = T883 ? io_in_bits_addr : inputReg_1_addr;
  assign T886 = inputReg_0_addr & T887;
  assign T887 = {6'h20/* 32*/{T888}};
  assign T888 = T6[1'h0/* 0*/];
  assign T889 = T843 && T890;
  assign T890 = T841[1'h0/* 0*/];
  assign T891 = T889 ? io_in_bits_addr : inputReg_0_addr;
  assign T892 = T896 && T893;
  assign T893 = ! T894;
  assign T894 = b == T895;
  assign T895 = {16'h0/* 0*/, 32'h6/* 6*/};
  assign T896 = T900 && T897;
  assign T897 = ! T898;
  assign T898 = b == T899;
  assign T899 = {16'h0/* 0*/, 32'h5/* 5*/};
  assign T900 = T904 && T901;
  assign T901 = ! T902;
  assign T902 = b == T903;
  assign T903 = {16'h0/* 0*/, 32'h4/* 4*/};
  assign T904 = T908 && T905;
  assign T905 = ! T906;
  assign T906 = b == T907;
  assign T907 = {16'h0/* 0*/, 32'h3/* 3*/};
  assign T908 = T912 && T909;
  assign T909 = ! T910;
  assign T910 = b == T911;
  assign T911 = {16'h0/* 0*/, 32'h2/* 2*/};
  assign T912 = T916 && T913;
  assign T913 = ! T914;
  assign T914 = b == T915;
  assign T915 = {16'h0/* 0*/, 32'h1/* 1*/};
  assign T916 = T920 && T917;
  assign T917 = ! T918;
  assign T918 = b == T919;
  assign T919 = {16'h0/* 0*/, 32'h0/* 0*/};
  assign T920 = T923 && T921;
  assign T921 = T768 == T922;
  assign T922 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T923 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T924 = T995 || T925;
  assign T925 = T926 && T777;
  assign T926 = T994 && T927;
  assign T927 = ! T928;
  assign T928 = T931 == r;
  assign r = T929 & 60'h7ffffff/* 134217727*/;
  assign T929 = {28'h0/* 0*/, T930};
  assign T930 = T836 >> 34'hf/* 15*/;
  assign T931 = {28'h0/* 0*/, T932};
  assign T932 = T940 | T933;
  assign T933 = rb7RowAddr_7 & T934;
  assign T934 = {6'h20/* 32*/{T5}};
  assign T935 = T839 || T936;
  assign T936 = T926 && T5;
  assign T937 = T936 ? r : T938;
  assign T938 = {28'h0/* 0*/, T939};
  assign T939 = T839 ? 32'h0/* 0*/ : rb7RowAddr_7;
  assign T940 = T948 | T941;
  assign T941 = rb7RowAddr_6 & T942;
  assign T942 = {6'h20/* 32*/{T764}};
  assign T943 = T849 || T944;
  assign T944 = T926 && T764;
  assign T945 = T944 ? r : T946;
  assign T946 = {28'h0/* 0*/, T947};
  assign T947 = T849 ? 32'h0/* 0*/ : rb7RowAddr_6;
  assign T948 = T955 | T949;
  assign T949 = rb7RowAddr_5 & T950;
  assign T950 = {6'h20/* 32*/{T777}};
  assign T951 = T855 || T925;
  assign T952 = T925 ? r : T953;
  assign T953 = {28'h0/* 0*/, T954};
  assign T954 = T855 ? 32'h0/* 0*/ : rb7RowAddr_5;
  assign T955 = T963 | T956;
  assign T956 = rb7RowAddr_4 & T957;
  assign T957 = {6'h20/* 32*/{T861}};
  assign T958 = T862 || T959;
  assign T959 = T926 && T861;
  assign T960 = T959 ? r : T961;
  assign T961 = {28'h0/* 0*/, T962};
  assign T962 = T862 ? 32'h0/* 0*/ : rb7RowAddr_4;
  assign T963 = T971 | T964;
  assign T964 = rb7RowAddr_3 & T965;
  assign T965 = {6'h20/* 32*/{T868}};
  assign T966 = T869 || T967;
  assign T967 = T926 && T868;
  assign T968 = T967 ? r : T969;
  assign T969 = {28'h0/* 0*/, T970};
  assign T970 = T869 ? 32'h0/* 0*/ : rb7RowAddr_3;
  assign T971 = T979 | T972;
  assign T972 = rb7RowAddr_2 & T973;
  assign T973 = {6'h20/* 32*/{T875}};
  assign T974 = T876 || T975;
  assign T975 = T926 && T875;
  assign T976 = T975 ? r : T977;
  assign T977 = {28'h0/* 0*/, T978};
  assign T978 = T876 ? 32'h0/* 0*/ : rb7RowAddr_2;
  assign T979 = T987 | T980;
  assign T980 = rb7RowAddr_1 & T981;
  assign T981 = {6'h20/* 32*/{T882}};
  assign T982 = T883 || T983;
  assign T983 = T926 && T882;
  assign T984 = T983 ? r : T985;
  assign T985 = {28'h0/* 0*/, T986};
  assign T986 = T883 ? 32'h0/* 0*/ : rb7RowAddr_1;
  assign T987 = rb7RowAddr_0 & T988;
  assign T988 = {6'h20/* 32*/{T888}};
  assign T989 = T889 || T990;
  assign T990 = T926 && T888;
  assign T991 = T990 ? r : T992;
  assign T992 = {28'h0/* 0*/, T993};
  assign T993 = T889 ? 32'h0/* 0*/ : rb7RowAddr_0;
  assign T994 = T892 && T832;
  assign T995 = T998 || T996;
  assign T996 = T997 && T777;
  assign T997 = T994 && T928;
  assign T998 = T1067 || T999;
  assign T999 = T1000 && T777;
  assign T1000 = T1066 && T1001;
  assign T1001 = ! T1002;
  assign T1002 = T1003 == r;
  assign T1003 = {28'h0/* 0*/, T1004};
  assign T1004 = T1012 | T1005;
  assign T1005 = rb6RowAddr_7 & T1006;
  assign T1006 = {6'h20/* 32*/{T5}};
  assign T1007 = T839 || T1008;
  assign T1008 = T1000 && T5;
  assign T1009 = T1008 ? r : T1010;
  assign T1010 = {28'h0/* 0*/, T1011};
  assign T1011 = T839 ? 32'h0/* 0*/ : rb6RowAddr_7;
  assign T1012 = T1020 | T1013;
  assign T1013 = rb6RowAddr_6 & T1014;
  assign T1014 = {6'h20/* 32*/{T764}};
  assign T1015 = T849 || T1016;
  assign T1016 = T1000 && T764;
  assign T1017 = T1016 ? r : T1018;
  assign T1018 = {28'h0/* 0*/, T1019};
  assign T1019 = T849 ? 32'h0/* 0*/ : rb6RowAddr_6;
  assign T1020 = T1027 | T1021;
  assign T1021 = rb6RowAddr_5 & T1022;
  assign T1022 = {6'h20/* 32*/{T777}};
  assign T1023 = T855 || T999;
  assign T1024 = T999 ? r : T1025;
  assign T1025 = {28'h0/* 0*/, T1026};
  assign T1026 = T855 ? 32'h0/* 0*/ : rb6RowAddr_5;
  assign T1027 = T1035 | T1028;
  assign T1028 = rb6RowAddr_4 & T1029;
  assign T1029 = {6'h20/* 32*/{T861}};
  assign T1030 = T862 || T1031;
  assign T1031 = T1000 && T861;
  assign T1032 = T1031 ? r : T1033;
  assign T1033 = {28'h0/* 0*/, T1034};
  assign T1034 = T862 ? 32'h0/* 0*/ : rb6RowAddr_4;
  assign T1035 = T1043 | T1036;
  assign T1036 = rb6RowAddr_3 & T1037;
  assign T1037 = {6'h20/* 32*/{T868}};
  assign T1038 = T869 || T1039;
  assign T1039 = T1000 && T868;
  assign T1040 = T1039 ? r : T1041;
  assign T1041 = {28'h0/* 0*/, T1042};
  assign T1042 = T869 ? 32'h0/* 0*/ : rb6RowAddr_3;
  assign T1043 = T1051 | T1044;
  assign T1044 = rb6RowAddr_2 & T1045;
  assign T1045 = {6'h20/* 32*/{T875}};
  assign T1046 = T876 || T1047;
  assign T1047 = T1000 && T875;
  assign T1048 = T1047 ? r : T1049;
  assign T1049 = {28'h0/* 0*/, T1050};
  assign T1050 = T876 ? 32'h0/* 0*/ : rb6RowAddr_2;
  assign T1051 = T1059 | T1052;
  assign T1052 = rb6RowAddr_1 & T1053;
  assign T1053 = {6'h20/* 32*/{T882}};
  assign T1054 = T883 || T1055;
  assign T1055 = T1000 && T882;
  assign T1056 = T1055 ? r : T1057;
  assign T1057 = {28'h0/* 0*/, T1058};
  assign T1058 = T883 ? 32'h0/* 0*/ : rb6RowAddr_1;
  assign T1059 = rb6RowAddr_0 & T1060;
  assign T1060 = {6'h20/* 32*/{T888}};
  assign T1061 = T889 || T1062;
  assign T1062 = T1000 && T888;
  assign T1063 = T1062 ? r : T1064;
  assign T1064 = {28'h0/* 0*/, T1065};
  assign T1065 = T889 ? 32'h0/* 0*/ : rb6RowAddr_0;
  assign T1066 = T896 && T894;
  assign T1067 = T1070 || T1068;
  assign T1068 = T1069 && T777;
  assign T1069 = T1066 && T1002;
  assign T1070 = T1139 || T1071;
  assign T1071 = T1072 && T777;
  assign T1072 = T1138 && T1073;
  assign T1073 = ! T1074;
  assign T1074 = T1075 == r;
  assign T1075 = {28'h0/* 0*/, T1076};
  assign T1076 = T1084 | T1077;
  assign T1077 = rb5RowAddr_7 & T1078;
  assign T1078 = {6'h20/* 32*/{T5}};
  assign T1079 = T839 || T1080;
  assign T1080 = T1072 && T5;
  assign T1081 = T1080 ? r : T1082;
  assign T1082 = {28'h0/* 0*/, T1083};
  assign T1083 = T839 ? 32'h0/* 0*/ : rb5RowAddr_7;
  assign T1084 = T1092 | T1085;
  assign T1085 = rb5RowAddr_6 & T1086;
  assign T1086 = {6'h20/* 32*/{T764}};
  assign T1087 = T849 || T1088;
  assign T1088 = T1072 && T764;
  assign T1089 = T1088 ? r : T1090;
  assign T1090 = {28'h0/* 0*/, T1091};
  assign T1091 = T849 ? 32'h0/* 0*/ : rb5RowAddr_6;
  assign T1092 = T1099 | T1093;
  assign T1093 = rb5RowAddr_5 & T1094;
  assign T1094 = {6'h20/* 32*/{T777}};
  assign T1095 = T855 || T1071;
  assign T1096 = T1071 ? r : T1097;
  assign T1097 = {28'h0/* 0*/, T1098};
  assign T1098 = T855 ? 32'h0/* 0*/ : rb5RowAddr_5;
  assign T1099 = T1107 | T1100;
  assign T1100 = rb5RowAddr_4 & T1101;
  assign T1101 = {6'h20/* 32*/{T861}};
  assign T1102 = T862 || T1103;
  assign T1103 = T1072 && T861;
  assign T1104 = T1103 ? r : T1105;
  assign T1105 = {28'h0/* 0*/, T1106};
  assign T1106 = T862 ? 32'h0/* 0*/ : rb5RowAddr_4;
  assign T1107 = T1115 | T1108;
  assign T1108 = rb5RowAddr_3 & T1109;
  assign T1109 = {6'h20/* 32*/{T868}};
  assign T1110 = T869 || T1111;
  assign T1111 = T1072 && T868;
  assign T1112 = T1111 ? r : T1113;
  assign T1113 = {28'h0/* 0*/, T1114};
  assign T1114 = T869 ? 32'h0/* 0*/ : rb5RowAddr_3;
  assign T1115 = T1123 | T1116;
  assign T1116 = rb5RowAddr_2 & T1117;
  assign T1117 = {6'h20/* 32*/{T875}};
  assign T1118 = T876 || T1119;
  assign T1119 = T1072 && T875;
  assign T1120 = T1119 ? r : T1121;
  assign T1121 = {28'h0/* 0*/, T1122};
  assign T1122 = T876 ? 32'h0/* 0*/ : rb5RowAddr_2;
  assign T1123 = T1131 | T1124;
  assign T1124 = rb5RowAddr_1 & T1125;
  assign T1125 = {6'h20/* 32*/{T882}};
  assign T1126 = T883 || T1127;
  assign T1127 = T1072 && T882;
  assign T1128 = T1127 ? r : T1129;
  assign T1129 = {28'h0/* 0*/, T1130};
  assign T1130 = T883 ? 32'h0/* 0*/ : rb5RowAddr_1;
  assign T1131 = rb5RowAddr_0 & T1132;
  assign T1132 = {6'h20/* 32*/{T888}};
  assign T1133 = T889 || T1134;
  assign T1134 = T1072 && T888;
  assign T1135 = T1134 ? r : T1136;
  assign T1136 = {28'h0/* 0*/, T1137};
  assign T1137 = T889 ? 32'h0/* 0*/ : rb5RowAddr_0;
  assign T1138 = T900 && T898;
  assign T1139 = T1142 || T1140;
  assign T1140 = T1141 && T777;
  assign T1141 = T1138 && T1074;
  assign T1142 = T1211 || T1143;
  assign T1143 = T1144 && T777;
  assign T1144 = T1210 && T1145;
  assign T1145 = ! T1146;
  assign T1146 = T1147 == r;
  assign T1147 = {28'h0/* 0*/, T1148};
  assign T1148 = T1156 | T1149;
  assign T1149 = rb4RowAddr_7 & T1150;
  assign T1150 = {6'h20/* 32*/{T5}};
  assign T1151 = T839 || T1152;
  assign T1152 = T1144 && T5;
  assign T1153 = T1152 ? r : T1154;
  assign T1154 = {28'h0/* 0*/, T1155};
  assign T1155 = T839 ? 32'h0/* 0*/ : rb4RowAddr_7;
  assign T1156 = T1164 | T1157;
  assign T1157 = rb4RowAddr_6 & T1158;
  assign T1158 = {6'h20/* 32*/{T764}};
  assign T1159 = T849 || T1160;
  assign T1160 = T1144 && T764;
  assign T1161 = T1160 ? r : T1162;
  assign T1162 = {28'h0/* 0*/, T1163};
  assign T1163 = T849 ? 32'h0/* 0*/ : rb4RowAddr_6;
  assign T1164 = T1171 | T1165;
  assign T1165 = rb4RowAddr_5 & T1166;
  assign T1166 = {6'h20/* 32*/{T777}};
  assign T1167 = T855 || T1143;
  assign T1168 = T1143 ? r : T1169;
  assign T1169 = {28'h0/* 0*/, T1170};
  assign T1170 = T855 ? 32'h0/* 0*/ : rb4RowAddr_5;
  assign T1171 = T1179 | T1172;
  assign T1172 = rb4RowAddr_4 & T1173;
  assign T1173 = {6'h20/* 32*/{T861}};
  assign T1174 = T862 || T1175;
  assign T1175 = T1144 && T861;
  assign T1176 = T1175 ? r : T1177;
  assign T1177 = {28'h0/* 0*/, T1178};
  assign T1178 = T862 ? 32'h0/* 0*/ : rb4RowAddr_4;
  assign T1179 = T1187 | T1180;
  assign T1180 = rb4RowAddr_3 & T1181;
  assign T1181 = {6'h20/* 32*/{T868}};
  assign T1182 = T869 || T1183;
  assign T1183 = T1144 && T868;
  assign T1184 = T1183 ? r : T1185;
  assign T1185 = {28'h0/* 0*/, T1186};
  assign T1186 = T869 ? 32'h0/* 0*/ : rb4RowAddr_3;
  assign T1187 = T1195 | T1188;
  assign T1188 = rb4RowAddr_2 & T1189;
  assign T1189 = {6'h20/* 32*/{T875}};
  assign T1190 = T876 || T1191;
  assign T1191 = T1144 && T875;
  assign T1192 = T1191 ? r : T1193;
  assign T1193 = {28'h0/* 0*/, T1194};
  assign T1194 = T876 ? 32'h0/* 0*/ : rb4RowAddr_2;
  assign T1195 = T1203 | T1196;
  assign T1196 = rb4RowAddr_1 & T1197;
  assign T1197 = {6'h20/* 32*/{T882}};
  assign T1198 = T883 || T1199;
  assign T1199 = T1144 && T882;
  assign T1200 = T1199 ? r : T1201;
  assign T1201 = {28'h0/* 0*/, T1202};
  assign T1202 = T883 ? 32'h0/* 0*/ : rb4RowAddr_1;
  assign T1203 = rb4RowAddr_0 & T1204;
  assign T1204 = {6'h20/* 32*/{T888}};
  assign T1205 = T889 || T1206;
  assign T1206 = T1144 && T888;
  assign T1207 = T1206 ? r : T1208;
  assign T1208 = {28'h0/* 0*/, T1209};
  assign T1209 = T889 ? 32'h0/* 0*/ : rb4RowAddr_0;
  assign T1210 = T904 && T902;
  assign T1211 = T1214 || T1212;
  assign T1212 = T1213 && T777;
  assign T1213 = T1210 && T1146;
  assign T1214 = T1283 || T1215;
  assign T1215 = T1216 && T777;
  assign T1216 = T1282 && T1217;
  assign T1217 = ! T1218;
  assign T1218 = T1219 == r;
  assign T1219 = {28'h0/* 0*/, T1220};
  assign T1220 = T1228 | T1221;
  assign T1221 = rb3RowAddr_7 & T1222;
  assign T1222 = {6'h20/* 32*/{T5}};
  assign T1223 = T839 || T1224;
  assign T1224 = T1216 && T5;
  assign T1225 = T1224 ? r : T1226;
  assign T1226 = {28'h0/* 0*/, T1227};
  assign T1227 = T839 ? 32'h0/* 0*/ : rb3RowAddr_7;
  assign T1228 = T1236 | T1229;
  assign T1229 = rb3RowAddr_6 & T1230;
  assign T1230 = {6'h20/* 32*/{T764}};
  assign T1231 = T849 || T1232;
  assign T1232 = T1216 && T764;
  assign T1233 = T1232 ? r : T1234;
  assign T1234 = {28'h0/* 0*/, T1235};
  assign T1235 = T849 ? 32'h0/* 0*/ : rb3RowAddr_6;
  assign T1236 = T1243 | T1237;
  assign T1237 = rb3RowAddr_5 & T1238;
  assign T1238 = {6'h20/* 32*/{T777}};
  assign T1239 = T855 || T1215;
  assign T1240 = T1215 ? r : T1241;
  assign T1241 = {28'h0/* 0*/, T1242};
  assign T1242 = T855 ? 32'h0/* 0*/ : rb3RowAddr_5;
  assign T1243 = T1251 | T1244;
  assign T1244 = rb3RowAddr_4 & T1245;
  assign T1245 = {6'h20/* 32*/{T861}};
  assign T1246 = T862 || T1247;
  assign T1247 = T1216 && T861;
  assign T1248 = T1247 ? r : T1249;
  assign T1249 = {28'h0/* 0*/, T1250};
  assign T1250 = T862 ? 32'h0/* 0*/ : rb3RowAddr_4;
  assign T1251 = T1259 | T1252;
  assign T1252 = rb3RowAddr_3 & T1253;
  assign T1253 = {6'h20/* 32*/{T868}};
  assign T1254 = T869 || T1255;
  assign T1255 = T1216 && T868;
  assign T1256 = T1255 ? r : T1257;
  assign T1257 = {28'h0/* 0*/, T1258};
  assign T1258 = T869 ? 32'h0/* 0*/ : rb3RowAddr_3;
  assign T1259 = T1267 | T1260;
  assign T1260 = rb3RowAddr_2 & T1261;
  assign T1261 = {6'h20/* 32*/{T875}};
  assign T1262 = T876 || T1263;
  assign T1263 = T1216 && T875;
  assign T1264 = T1263 ? r : T1265;
  assign T1265 = {28'h0/* 0*/, T1266};
  assign T1266 = T876 ? 32'h0/* 0*/ : rb3RowAddr_2;
  assign T1267 = T1275 | T1268;
  assign T1268 = rb3RowAddr_1 & T1269;
  assign T1269 = {6'h20/* 32*/{T882}};
  assign T1270 = T883 || T1271;
  assign T1271 = T1216 && T882;
  assign T1272 = T1271 ? r : T1273;
  assign T1273 = {28'h0/* 0*/, T1274};
  assign T1274 = T883 ? 32'h0/* 0*/ : rb3RowAddr_1;
  assign T1275 = rb3RowAddr_0 & T1276;
  assign T1276 = {6'h20/* 32*/{T888}};
  assign T1277 = T889 || T1278;
  assign T1278 = T1216 && T888;
  assign T1279 = T1278 ? r : T1280;
  assign T1280 = {28'h0/* 0*/, T1281};
  assign T1281 = T889 ? 32'h0/* 0*/ : rb3RowAddr_0;
  assign T1282 = T908 && T906;
  assign T1283 = T1286 || T1284;
  assign T1284 = T1285 && T777;
  assign T1285 = T1282 && T1218;
  assign T1286 = T1355 || T1287;
  assign T1287 = T1288 && T777;
  assign T1288 = T1354 && T1289;
  assign T1289 = ! T1290;
  assign T1290 = T1291 == r;
  assign T1291 = {28'h0/* 0*/, T1292};
  assign T1292 = T1300 | T1293;
  assign T1293 = rb2RowAddr_7 & T1294;
  assign T1294 = {6'h20/* 32*/{T5}};
  assign T1295 = T839 || T1296;
  assign T1296 = T1288 && T5;
  assign T1297 = T1296 ? r : T1298;
  assign T1298 = {28'h0/* 0*/, T1299};
  assign T1299 = T839 ? 32'h0/* 0*/ : rb2RowAddr_7;
  assign T1300 = T1308 | T1301;
  assign T1301 = rb2RowAddr_6 & T1302;
  assign T1302 = {6'h20/* 32*/{T764}};
  assign T1303 = T849 || T1304;
  assign T1304 = T1288 && T764;
  assign T1305 = T1304 ? r : T1306;
  assign T1306 = {28'h0/* 0*/, T1307};
  assign T1307 = T849 ? 32'h0/* 0*/ : rb2RowAddr_6;
  assign T1308 = T1315 | T1309;
  assign T1309 = rb2RowAddr_5 & T1310;
  assign T1310 = {6'h20/* 32*/{T777}};
  assign T1311 = T855 || T1287;
  assign T1312 = T1287 ? r : T1313;
  assign T1313 = {28'h0/* 0*/, T1314};
  assign T1314 = T855 ? 32'h0/* 0*/ : rb2RowAddr_5;
  assign T1315 = T1323 | T1316;
  assign T1316 = rb2RowAddr_4 & T1317;
  assign T1317 = {6'h20/* 32*/{T861}};
  assign T1318 = T862 || T1319;
  assign T1319 = T1288 && T861;
  assign T1320 = T1319 ? r : T1321;
  assign T1321 = {28'h0/* 0*/, T1322};
  assign T1322 = T862 ? 32'h0/* 0*/ : rb2RowAddr_4;
  assign T1323 = T1331 | T1324;
  assign T1324 = rb2RowAddr_3 & T1325;
  assign T1325 = {6'h20/* 32*/{T868}};
  assign T1326 = T869 || T1327;
  assign T1327 = T1288 && T868;
  assign T1328 = T1327 ? r : T1329;
  assign T1329 = {28'h0/* 0*/, T1330};
  assign T1330 = T869 ? 32'h0/* 0*/ : rb2RowAddr_3;
  assign T1331 = T1339 | T1332;
  assign T1332 = rb2RowAddr_2 & T1333;
  assign T1333 = {6'h20/* 32*/{T875}};
  assign T1334 = T876 || T1335;
  assign T1335 = T1288 && T875;
  assign T1336 = T1335 ? r : T1337;
  assign T1337 = {28'h0/* 0*/, T1338};
  assign T1338 = T876 ? 32'h0/* 0*/ : rb2RowAddr_2;
  assign T1339 = T1347 | T1340;
  assign T1340 = rb2RowAddr_1 & T1341;
  assign T1341 = {6'h20/* 32*/{T882}};
  assign T1342 = T883 || T1343;
  assign T1343 = T1288 && T882;
  assign T1344 = T1343 ? r : T1345;
  assign T1345 = {28'h0/* 0*/, T1346};
  assign T1346 = T883 ? 32'h0/* 0*/ : rb2RowAddr_1;
  assign T1347 = rb2RowAddr_0 & T1348;
  assign T1348 = {6'h20/* 32*/{T888}};
  assign T1349 = T889 || T1350;
  assign T1350 = T1288 && T888;
  assign T1351 = T1350 ? r : T1352;
  assign T1352 = {28'h0/* 0*/, T1353};
  assign T1353 = T889 ? 32'h0/* 0*/ : rb2RowAddr_0;
  assign T1354 = T912 && T910;
  assign T1355 = T1358 || T1356;
  assign T1356 = T1357 && T777;
  assign T1357 = T1354 && T1290;
  assign T1358 = T1427 || T1359;
  assign T1359 = T1360 && T777;
  assign T1360 = T1426 && T1361;
  assign T1361 = ! T1362;
  assign T1362 = T1363 == r;
  assign T1363 = {28'h0/* 0*/, T1364};
  assign T1364 = T1372 | T1365;
  assign T1365 = rb1RowAddr_7 & T1366;
  assign T1366 = {6'h20/* 32*/{T5}};
  assign T1367 = T839 || T1368;
  assign T1368 = T1360 && T5;
  assign T1369 = T1368 ? r : T1370;
  assign T1370 = {28'h0/* 0*/, T1371};
  assign T1371 = T839 ? 32'h0/* 0*/ : rb1RowAddr_7;
  assign T1372 = T1380 | T1373;
  assign T1373 = rb1RowAddr_6 & T1374;
  assign T1374 = {6'h20/* 32*/{T764}};
  assign T1375 = T849 || T1376;
  assign T1376 = T1360 && T764;
  assign T1377 = T1376 ? r : T1378;
  assign T1378 = {28'h0/* 0*/, T1379};
  assign T1379 = T849 ? 32'h0/* 0*/ : rb1RowAddr_6;
  assign T1380 = T1387 | T1381;
  assign T1381 = rb1RowAddr_5 & T1382;
  assign T1382 = {6'h20/* 32*/{T777}};
  assign T1383 = T855 || T1359;
  assign T1384 = T1359 ? r : T1385;
  assign T1385 = {28'h0/* 0*/, T1386};
  assign T1386 = T855 ? 32'h0/* 0*/ : rb1RowAddr_5;
  assign T1387 = T1395 | T1388;
  assign T1388 = rb1RowAddr_4 & T1389;
  assign T1389 = {6'h20/* 32*/{T861}};
  assign T1390 = T862 || T1391;
  assign T1391 = T1360 && T861;
  assign T1392 = T1391 ? r : T1393;
  assign T1393 = {28'h0/* 0*/, T1394};
  assign T1394 = T862 ? 32'h0/* 0*/ : rb1RowAddr_4;
  assign T1395 = T1403 | T1396;
  assign T1396 = rb1RowAddr_3 & T1397;
  assign T1397 = {6'h20/* 32*/{T868}};
  assign T1398 = T869 || T1399;
  assign T1399 = T1360 && T868;
  assign T1400 = T1399 ? r : T1401;
  assign T1401 = {28'h0/* 0*/, T1402};
  assign T1402 = T869 ? 32'h0/* 0*/ : rb1RowAddr_3;
  assign T1403 = T1411 | T1404;
  assign T1404 = rb1RowAddr_2 & T1405;
  assign T1405 = {6'h20/* 32*/{T875}};
  assign T1406 = T876 || T1407;
  assign T1407 = T1360 && T875;
  assign T1408 = T1407 ? r : T1409;
  assign T1409 = {28'h0/* 0*/, T1410};
  assign T1410 = T876 ? 32'h0/* 0*/ : rb1RowAddr_2;
  assign T1411 = T1419 | T1412;
  assign T1412 = rb1RowAddr_1 & T1413;
  assign T1413 = {6'h20/* 32*/{T882}};
  assign T1414 = T883 || T1415;
  assign T1415 = T1360 && T882;
  assign T1416 = T1415 ? r : T1417;
  assign T1417 = {28'h0/* 0*/, T1418};
  assign T1418 = T883 ? 32'h0/* 0*/ : rb1RowAddr_1;
  assign T1419 = rb1RowAddr_0 & T1420;
  assign T1420 = {6'h20/* 32*/{T888}};
  assign T1421 = T889 || T1422;
  assign T1422 = T1360 && T888;
  assign T1423 = T1422 ? r : T1424;
  assign T1424 = {28'h0/* 0*/, T1425};
  assign T1425 = T889 ? 32'h0/* 0*/ : rb1RowAddr_0;
  assign T1426 = T916 && T914;
  assign T1427 = T1430 || T1428;
  assign T1428 = T1429 && T777;
  assign T1429 = T1426 && T1362;
  assign T1430 = T1499 || T1431;
  assign T1431 = T1432 && T777;
  assign T1432 = T1498 && T1433;
  assign T1433 = ! T1434;
  assign T1434 = T1435 == r;
  assign T1435 = {28'h0/* 0*/, T1436};
  assign T1436 = T1444 | T1437;
  assign T1437 = rb0RowAddr_7 & T1438;
  assign T1438 = {6'h20/* 32*/{T5}};
  assign T1439 = T839 || T1440;
  assign T1440 = T1432 && T5;
  assign T1441 = T1440 ? r : T1442;
  assign T1442 = {28'h0/* 0*/, T1443};
  assign T1443 = T839 ? 32'h1/* 1*/ : rb0RowAddr_7;
  assign T1444 = T1452 | T1445;
  assign T1445 = rb0RowAddr_6 & T1446;
  assign T1446 = {6'h20/* 32*/{T764}};
  assign T1447 = T849 || T1448;
  assign T1448 = T1432 && T764;
  assign T1449 = T1448 ? r : T1450;
  assign T1450 = {28'h0/* 0*/, T1451};
  assign T1451 = T849 ? 32'h1/* 1*/ : rb0RowAddr_6;
  assign T1452 = T1459 | T1453;
  assign T1453 = rb0RowAddr_5 & T1454;
  assign T1454 = {6'h20/* 32*/{T777}};
  assign T1455 = T855 || T1431;
  assign T1456 = T1431 ? r : T1457;
  assign T1457 = {28'h0/* 0*/, T1458};
  assign T1458 = T855 ? 32'h1/* 1*/ : rb0RowAddr_5;
  assign T1459 = T1467 | T1460;
  assign T1460 = rb0RowAddr_4 & T1461;
  assign T1461 = {6'h20/* 32*/{T861}};
  assign T1462 = T862 || T1463;
  assign T1463 = T1432 && T861;
  assign T1464 = T1463 ? r : T1465;
  assign T1465 = {28'h0/* 0*/, T1466};
  assign T1466 = T862 ? 32'h1/* 1*/ : rb0RowAddr_4;
  assign T1467 = T1475 | T1468;
  assign T1468 = rb0RowAddr_3 & T1469;
  assign T1469 = {6'h20/* 32*/{T868}};
  assign T1470 = T869 || T1471;
  assign T1471 = T1432 && T868;
  assign T1472 = T1471 ? r : T1473;
  assign T1473 = {28'h0/* 0*/, T1474};
  assign T1474 = T869 ? 32'h1/* 1*/ : rb0RowAddr_3;
  assign T1475 = T1483 | T1476;
  assign T1476 = rb0RowAddr_2 & T1477;
  assign T1477 = {6'h20/* 32*/{T875}};
  assign T1478 = T876 || T1479;
  assign T1479 = T1432 && T875;
  assign T1480 = T1479 ? r : T1481;
  assign T1481 = {28'h0/* 0*/, T1482};
  assign T1482 = T876 ? 32'h1/* 1*/ : rb0RowAddr_2;
  assign T1483 = T1491 | T1484;
  assign T1484 = rb0RowAddr_1 & T1485;
  assign T1485 = {6'h20/* 32*/{T882}};
  assign T1486 = T883 || T1487;
  assign T1487 = T1432 && T882;
  assign T1488 = T1487 ? r : T1489;
  assign T1489 = {28'h0/* 0*/, T1490};
  assign T1490 = T883 ? 32'h1/* 1*/ : rb0RowAddr_1;
  assign T1491 = rb0RowAddr_0 & T1492;
  assign T1492 = {6'h20/* 32*/{T888}};
  assign T1493 = T889 || T1494;
  assign T1494 = T1432 && T888;
  assign T1495 = T1494 ? r : T1496;
  assign T1496 = {28'h0/* 0*/, T1497};
  assign T1497 = T889 ? 32'h1/* 1*/ : rb0RowAddr_0;
  assign T1498 = T920 && T918;
  assign T1499 = T1502 || T1500;
  assign T1500 = T1501 && T777;
  assign T1501 = T1498 && T1434;
  assign T1502 = T855 || T1503;
  assign T1503 = T1504 && T84;
  assign T1504 = T1505 && io_out_ready;
  assign T1505 = T1507 && T1506;
  assign T1506 = T19 == 8'hff/* 255*/;
  assign T1507 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T1508 = T1766 ? 8'hff/* 255*/ : T1509;
  assign T1509 = T829 ? T1765 : T1510;
  assign T1510 = T925 ? T1764 : T1511;
  assign T1511 = T996 ? T1763 : T1512;
  assign T1512 = T999 ? T1762 : T1513;
  assign T1513 = T1068 ? T1761 : T1514;
  assign T1514 = T1071 ? T1760 : T1515;
  assign T1515 = T1140 ? T1759 : T1516;
  assign T1516 = T1143 ? T1758 : T1517;
  assign T1517 = T1212 ? T1757 : T1518;
  assign T1518 = T1215 ? T1756 : T1519;
  assign T1519 = T1284 ? T1755 : T1520;
  assign T1520 = T1287 ? T1754 : T1521;
  assign T1521 = T1356 ? T1753 : T1522;
  assign T1522 = T1359 ? T1752 : T1523;
  assign T1523 = T1428 ? T1751 : T1524;
  assign T1524 = T1431 ? T1750 : T1525;
  assign T1525 = T1500 ? T1749 : T1526;
  assign T1526 = T1503 ? T1529 : T1527;
  assign T1527 = T855 ? T1528 : State_5;
  assign T1528 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1529 = T1557 | T1530;
  assign T1530 = EmitReturnState_7 & T1531;
  assign T1531 = {4'h8/* 8*/{T22}};
  assign T1532 = T1533 || T4;
  assign T1533 = T1535 || T1534;
  assign T1534 = T782 && T5;
  assign T1535 = T1537 || T1536;
  assign T1536 = T788 && T5;
  assign T1537 = T1539 || T1538;
  assign T1538 = T794 && T5;
  assign T1539 = T1541 || T1540;
  assign T1540 = T800 && T5;
  assign T1541 = T1543 || T1542;
  assign T1542 = T806 && T5;
  assign T1543 = T1545 || T1544;
  assign T1544 = T812 && T5;
  assign T1545 = T1547 || T1546;
  assign T1546 = T818 && T5;
  assign T1547 = T824 && T5;
  assign T1548 = T1549 ? 8'h0/* 0*/ : EmitReturnState_7;
  assign T1549 = T1550 || T4;
  assign T1550 = T1551 || T1534;
  assign T1551 = T1552 || T1536;
  assign T1552 = T1553 || T1538;
  assign T1553 = T1554 || T1540;
  assign T1554 = T1555 || T1542;
  assign T1555 = T1556 || T1544;
  assign T1556 = T1547 || T1546;
  assign T1557 = T1585 | T1558;
  assign T1558 = EmitReturnState_6 & T1559;
  assign T1559 = {4'h8/* 8*/{T73}};
  assign T1560 = T1561 || T763;
  assign T1561 = T1563 || T1562;
  assign T1562 = T782 && T764;
  assign T1563 = T1565 || T1564;
  assign T1564 = T788 && T764;
  assign T1565 = T1567 || T1566;
  assign T1566 = T794 && T764;
  assign T1567 = T1569 || T1568;
  assign T1568 = T800 && T764;
  assign T1569 = T1571 || T1570;
  assign T1570 = T806 && T764;
  assign T1571 = T1573 || T1572;
  assign T1572 = T812 && T764;
  assign T1573 = T1575 || T1574;
  assign T1574 = T818 && T764;
  assign T1575 = T824 && T764;
  assign T1576 = T1577 ? 8'h0/* 0*/ : EmitReturnState_6;
  assign T1577 = T1578 || T763;
  assign T1578 = T1579 || T1562;
  assign T1579 = T1580 || T1564;
  assign T1580 = T1581 || T1566;
  assign T1581 = T1582 || T1568;
  assign T1582 = T1583 || T1570;
  assign T1583 = T1584 || T1572;
  assign T1584 = T1575 || T1574;
  assign T1585 = T1605 | T1586;
  assign T1586 = EmitReturnState_5 & T1587;
  assign T1587 = {4'h8/* 8*/{T84}};
  assign T1588 = T1589 || T779;
  assign T1589 = T1590 || T781;
  assign T1590 = T1591 || T787;
  assign T1591 = T1592 || T793;
  assign T1592 = T1593 || T799;
  assign T1593 = T1594 || T805;
  assign T1594 = T1595 || T811;
  assign T1595 = T823 || T817;
  assign T1596 = T1597 ? 8'h0/* 0*/ : EmitReturnState_5;
  assign T1597 = T1598 || T779;
  assign T1598 = T1599 || T781;
  assign T1599 = T1600 || T787;
  assign T1600 = T1601 || T793;
  assign T1601 = T1602 || T799;
  assign T1602 = T1603 || T805;
  assign T1603 = T1604 || T811;
  assign T1604 = T823 || T817;
  assign T1605 = T1634 | T1606;
  assign T1606 = EmitReturnState_4 & T1607;
  assign T1607 = {4'h8/* 8*/{T95}};
  assign T1608 = T1610 || T1609;
  assign T1609 = T765 && T861;
  assign T1610 = T1612 || T1611;
  assign T1611 = T782 && T861;
  assign T1612 = T1614 || T1613;
  assign T1613 = T788 && T861;
  assign T1614 = T1616 || T1615;
  assign T1615 = T794 && T861;
  assign T1616 = T1618 || T1617;
  assign T1617 = T800 && T861;
  assign T1618 = T1620 || T1619;
  assign T1619 = T806 && T861;
  assign T1620 = T1622 || T1621;
  assign T1621 = T812 && T861;
  assign T1622 = T1624 || T1623;
  assign T1623 = T818 && T861;
  assign T1624 = T824 && T861;
  assign T1625 = T1626 ? 8'h0/* 0*/ : EmitReturnState_4;
  assign T1626 = T1627 || T1609;
  assign T1627 = T1628 || T1611;
  assign T1628 = T1629 || T1613;
  assign T1629 = T1630 || T1615;
  assign T1630 = T1631 || T1617;
  assign T1631 = T1632 || T1619;
  assign T1632 = T1633 || T1621;
  assign T1633 = T1624 || T1623;
  assign T1634 = T1663 | T1635;
  assign T1635 = EmitReturnState_3 & T1636;
  assign T1636 = {4'h8/* 8*/{T106}};
  assign T1637 = T1639 || T1638;
  assign T1638 = T765 && T868;
  assign T1639 = T1641 || T1640;
  assign T1640 = T782 && T868;
  assign T1641 = T1643 || T1642;
  assign T1642 = T788 && T868;
  assign T1643 = T1645 || T1644;
  assign T1644 = T794 && T868;
  assign T1645 = T1647 || T1646;
  assign T1646 = T800 && T868;
  assign T1647 = T1649 || T1648;
  assign T1648 = T806 && T868;
  assign T1649 = T1651 || T1650;
  assign T1650 = T812 && T868;
  assign T1651 = T1653 || T1652;
  assign T1652 = T818 && T868;
  assign T1653 = T824 && T868;
  assign T1654 = T1655 ? 8'h0/* 0*/ : EmitReturnState_3;
  assign T1655 = T1656 || T1638;
  assign T1656 = T1657 || T1640;
  assign T1657 = T1658 || T1642;
  assign T1658 = T1659 || T1644;
  assign T1659 = T1660 || T1646;
  assign T1660 = T1661 || T1648;
  assign T1661 = T1662 || T1650;
  assign T1662 = T1653 || T1652;
  assign T1663 = T1692 | T1664;
  assign T1664 = EmitReturnState_2 & T1665;
  assign T1665 = {4'h8/* 8*/{T117}};
  assign T1666 = T1668 || T1667;
  assign T1667 = T765 && T875;
  assign T1668 = T1670 || T1669;
  assign T1669 = T782 && T875;
  assign T1670 = T1672 || T1671;
  assign T1671 = T788 && T875;
  assign T1672 = T1674 || T1673;
  assign T1673 = T794 && T875;
  assign T1674 = T1676 || T1675;
  assign T1675 = T800 && T875;
  assign T1676 = T1678 || T1677;
  assign T1677 = T806 && T875;
  assign T1678 = T1680 || T1679;
  assign T1679 = T812 && T875;
  assign T1680 = T1682 || T1681;
  assign T1681 = T818 && T875;
  assign T1682 = T824 && T875;
  assign T1683 = T1684 ? 8'h0/* 0*/ : EmitReturnState_2;
  assign T1684 = T1685 || T1667;
  assign T1685 = T1686 || T1669;
  assign T1686 = T1687 || T1671;
  assign T1687 = T1688 || T1673;
  assign T1688 = T1689 || T1675;
  assign T1689 = T1690 || T1677;
  assign T1690 = T1691 || T1679;
  assign T1691 = T1682 || T1681;
  assign T1692 = T1721 | T1693;
  assign T1693 = EmitReturnState_1 & T1694;
  assign T1694 = {4'h8/* 8*/{T128}};
  assign T1695 = T1697 || T1696;
  assign T1696 = T765 && T882;
  assign T1697 = T1699 || T1698;
  assign T1698 = T782 && T882;
  assign T1699 = T1701 || T1700;
  assign T1700 = T788 && T882;
  assign T1701 = T1703 || T1702;
  assign T1702 = T794 && T882;
  assign T1703 = T1705 || T1704;
  assign T1704 = T800 && T882;
  assign T1705 = T1707 || T1706;
  assign T1706 = T806 && T882;
  assign T1707 = T1709 || T1708;
  assign T1708 = T812 && T882;
  assign T1709 = T1711 || T1710;
  assign T1710 = T818 && T882;
  assign T1711 = T824 && T882;
  assign T1712 = T1713 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T1713 = T1714 || T1696;
  assign T1714 = T1715 || T1698;
  assign T1715 = T1716 || T1700;
  assign T1716 = T1717 || T1702;
  assign T1717 = T1718 || T1704;
  assign T1718 = T1719 || T1706;
  assign T1719 = T1720 || T1708;
  assign T1720 = T1711 || T1710;
  assign T1721 = EmitReturnState_0 & T1722;
  assign T1722 = {4'h8/* 8*/{T138}};
  assign T1723 = T1725 || T1724;
  assign T1724 = T765 && T888;
  assign T1725 = T1727 || T1726;
  assign T1726 = T782 && T888;
  assign T1727 = T1729 || T1728;
  assign T1728 = T788 && T888;
  assign T1729 = T1731 || T1730;
  assign T1730 = T794 && T888;
  assign T1731 = T1733 || T1732;
  assign T1732 = T800 && T888;
  assign T1733 = T1735 || T1734;
  assign T1734 = T806 && T888;
  assign T1735 = T1737 || T1736;
  assign T1736 = T812 && T888;
  assign T1737 = T1739 || T1738;
  assign T1738 = T818 && T888;
  assign T1739 = T824 && T888;
  assign T1740 = T1741 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T1741 = T1742 || T1724;
  assign T1742 = T1743 || T1726;
  assign T1743 = T1744 || T1728;
  assign T1744 = T1745 || T1730;
  assign T1745 = T1746 || T1732;
  assign T1746 = T1747 || T1734;
  assign T1747 = T1748 || T1736;
  assign T1748 = T1739 || T1738;
  assign T1749 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1750 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1751 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1752 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1753 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1754 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1755 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1756 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1757 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1758 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1759 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1760 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1761 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1762 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1763 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1764 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1765 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1766 = T1767 || T779;
  assign T1767 = T1768 || T781;
  assign T1768 = T1769 || T787;
  assign T1769 = T1770 || T793;
  assign T1770 = T1771 || T799;
  assign T1771 = T1772 || T805;
  assign T1772 = T1773 || T811;
  assign T1773 = T823 || T817;
  assign T1774 = T1860 | T1775;
  assign T1775 = State_4 & T1776;
  assign T1776 = {4'h8/* 8*/{T861}};
  assign T1777 = T1778 || T1609;
  assign T1778 = T1779 || T1611;
  assign T1779 = T1780 || T1613;
  assign T1780 = T1781 || T1615;
  assign T1781 = T1782 || T1617;
  assign T1782 = T1783 || T1619;
  assign T1783 = T1784 || T1621;
  assign T1784 = T1785 || T1623;
  assign T1785 = T1786 || T1624;
  assign T1786 = T1788 || T1787;
  assign T1787 = T830 && T861;
  assign T1788 = T1789 || T959;
  assign T1789 = T1791 || T1790;
  assign T1790 = T997 && T861;
  assign T1791 = T1792 || T1031;
  assign T1792 = T1794 || T1793;
  assign T1793 = T1069 && T861;
  assign T1794 = T1795 || T1103;
  assign T1795 = T1797 || T1796;
  assign T1796 = T1141 && T861;
  assign T1797 = T1798 || T1175;
  assign T1798 = T1800 || T1799;
  assign T1799 = T1213 && T861;
  assign T1800 = T1801 || T1247;
  assign T1801 = T1803 || T1802;
  assign T1802 = T1285 && T861;
  assign T1803 = T1804 || T1319;
  assign T1804 = T1806 || T1805;
  assign T1805 = T1357 && T861;
  assign T1806 = T1807 || T1391;
  assign T1807 = T1809 || T1808;
  assign T1808 = T1429 && T861;
  assign T1809 = T1810 || T1463;
  assign T1810 = T1812 || T1811;
  assign T1811 = T1501 && T861;
  assign T1812 = T862 || T1813;
  assign T1813 = T1504 && T95;
  assign T1814 = T1852 ? 8'hff/* 255*/ : T1815;
  assign T1815 = T1787 ? T1851 : T1816;
  assign T1816 = T959 ? T1850 : T1817;
  assign T1817 = T1790 ? T1849 : T1818;
  assign T1818 = T1031 ? T1848 : T1819;
  assign T1819 = T1793 ? T1847 : T1820;
  assign T1820 = T1103 ? T1846 : T1821;
  assign T1821 = T1796 ? T1845 : T1822;
  assign T1822 = T1175 ? T1844 : T1823;
  assign T1823 = T1799 ? T1843 : T1824;
  assign T1824 = T1247 ? T1842 : T1825;
  assign T1825 = T1802 ? T1841 : T1826;
  assign T1826 = T1319 ? T1840 : T1827;
  assign T1827 = T1805 ? T1839 : T1828;
  assign T1828 = T1391 ? T1838 : T1829;
  assign T1829 = T1808 ? T1837 : T1830;
  assign T1830 = T1463 ? T1836 : T1831;
  assign T1831 = T1811 ? T1835 : T1832;
  assign T1832 = T1813 ? T1529 : T1833;
  assign T1833 = T862 ? T1834 : State_4;
  assign T1834 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1835 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1836 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1837 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1838 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1839 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1840 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1841 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1842 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1843 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1844 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1845 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1846 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1847 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1848 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1849 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1850 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1851 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1852 = T1853 || T1609;
  assign T1853 = T1854 || T1611;
  assign T1854 = T1855 || T1613;
  assign T1855 = T1856 || T1615;
  assign T1856 = T1857 || T1617;
  assign T1857 = T1858 || T1619;
  assign T1858 = T1859 || T1621;
  assign T1859 = T1624 || T1623;
  assign T1860 = T1946 | T1861;
  assign T1861 = State_3 & T1862;
  assign T1862 = {4'h8/* 8*/{T868}};
  assign T1863 = T1864 || T1638;
  assign T1864 = T1865 || T1640;
  assign T1865 = T1866 || T1642;
  assign T1866 = T1867 || T1644;
  assign T1867 = T1868 || T1646;
  assign T1868 = T1869 || T1648;
  assign T1869 = T1870 || T1650;
  assign T1870 = T1871 || T1652;
  assign T1871 = T1872 || T1653;
  assign T1872 = T1874 || T1873;
  assign T1873 = T830 && T868;
  assign T1874 = T1875 || T967;
  assign T1875 = T1877 || T1876;
  assign T1876 = T997 && T868;
  assign T1877 = T1878 || T1039;
  assign T1878 = T1880 || T1879;
  assign T1879 = T1069 && T868;
  assign T1880 = T1881 || T1111;
  assign T1881 = T1883 || T1882;
  assign T1882 = T1141 && T868;
  assign T1883 = T1884 || T1183;
  assign T1884 = T1886 || T1885;
  assign T1885 = T1213 && T868;
  assign T1886 = T1887 || T1255;
  assign T1887 = T1889 || T1888;
  assign T1888 = T1285 && T868;
  assign T1889 = T1890 || T1327;
  assign T1890 = T1892 || T1891;
  assign T1891 = T1357 && T868;
  assign T1892 = T1893 || T1399;
  assign T1893 = T1895 || T1894;
  assign T1894 = T1429 && T868;
  assign T1895 = T1896 || T1471;
  assign T1896 = T1898 || T1897;
  assign T1897 = T1501 && T868;
  assign T1898 = T869 || T1899;
  assign T1899 = T1504 && T106;
  assign T1900 = T1938 ? 8'hff/* 255*/ : T1901;
  assign T1901 = T1873 ? T1937 : T1902;
  assign T1902 = T967 ? T1936 : T1903;
  assign T1903 = T1876 ? T1935 : T1904;
  assign T1904 = T1039 ? T1934 : T1905;
  assign T1905 = T1879 ? T1933 : T1906;
  assign T1906 = T1111 ? T1932 : T1907;
  assign T1907 = T1882 ? T1931 : T1908;
  assign T1908 = T1183 ? T1930 : T1909;
  assign T1909 = T1885 ? T1929 : T1910;
  assign T1910 = T1255 ? T1928 : T1911;
  assign T1911 = T1888 ? T1927 : T1912;
  assign T1912 = T1327 ? T1926 : T1913;
  assign T1913 = T1891 ? T1925 : T1914;
  assign T1914 = T1399 ? T1924 : T1915;
  assign T1915 = T1894 ? T1923 : T1916;
  assign T1916 = T1471 ? T1922 : T1917;
  assign T1917 = T1897 ? T1921 : T1918;
  assign T1918 = T1899 ? T1529 : T1919;
  assign T1919 = T869 ? T1920 : State_3;
  assign T1920 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1921 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1922 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1923 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1924 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1925 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1926 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1927 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1928 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1929 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1930 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1931 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1932 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1933 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1934 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1935 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1936 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1937 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1938 = T1939 || T1638;
  assign T1939 = T1940 || T1640;
  assign T1940 = T1941 || T1642;
  assign T1941 = T1942 || T1644;
  assign T1942 = T1943 || T1646;
  assign T1943 = T1944 || T1648;
  assign T1944 = T1945 || T1650;
  assign T1945 = T1653 || T1652;
  assign T1946 = T2032 | T1947;
  assign T1947 = State_2 & T1948;
  assign T1948 = {4'h8/* 8*/{T875}};
  assign T1949 = T1950 || T1667;
  assign T1950 = T1951 || T1669;
  assign T1951 = T1952 || T1671;
  assign T1952 = T1953 || T1673;
  assign T1953 = T1954 || T1675;
  assign T1954 = T1955 || T1677;
  assign T1955 = T1956 || T1679;
  assign T1956 = T1957 || T1681;
  assign T1957 = T1958 || T1682;
  assign T1958 = T1960 || T1959;
  assign T1959 = T830 && T875;
  assign T1960 = T1961 || T975;
  assign T1961 = T1963 || T1962;
  assign T1962 = T997 && T875;
  assign T1963 = T1964 || T1047;
  assign T1964 = T1966 || T1965;
  assign T1965 = T1069 && T875;
  assign T1966 = T1967 || T1119;
  assign T1967 = T1969 || T1968;
  assign T1968 = T1141 && T875;
  assign T1969 = T1970 || T1191;
  assign T1970 = T1972 || T1971;
  assign T1971 = T1213 && T875;
  assign T1972 = T1973 || T1263;
  assign T1973 = T1975 || T1974;
  assign T1974 = T1285 && T875;
  assign T1975 = T1976 || T1335;
  assign T1976 = T1978 || T1977;
  assign T1977 = T1357 && T875;
  assign T1978 = T1979 || T1407;
  assign T1979 = T1981 || T1980;
  assign T1980 = T1429 && T875;
  assign T1981 = T1982 || T1479;
  assign T1982 = T1984 || T1983;
  assign T1983 = T1501 && T875;
  assign T1984 = T876 || T1985;
  assign T1985 = T1504 && T117;
  assign T1986 = T2024 ? 8'hff/* 255*/ : T1987;
  assign T1987 = T1959 ? T2023 : T1988;
  assign T1988 = T975 ? T2022 : T1989;
  assign T1989 = T1962 ? T2021 : T1990;
  assign T1990 = T1047 ? T2020 : T1991;
  assign T1991 = T1965 ? T2019 : T1992;
  assign T1992 = T1119 ? T2018 : T1993;
  assign T1993 = T1968 ? T2017 : T1994;
  assign T1994 = T1191 ? T2016 : T1995;
  assign T1995 = T1971 ? T2015 : T1996;
  assign T1996 = T1263 ? T2014 : T1997;
  assign T1997 = T1974 ? T2013 : T1998;
  assign T1998 = T1335 ? T2012 : T1999;
  assign T1999 = T1977 ? T2011 : T2000;
  assign T2000 = T1407 ? T2010 : T2001;
  assign T2001 = T1980 ? T2009 : T2002;
  assign T2002 = T1479 ? T2008 : T2003;
  assign T2003 = T1983 ? T2007 : T2004;
  assign T2004 = T1985 ? T1529 : T2005;
  assign T2005 = T876 ? T2006 : State_2;
  assign T2006 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2007 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2008 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2009 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2010 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2011 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2012 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2013 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2014 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2015 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2016 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2017 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2018 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2019 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2020 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2021 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2022 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2023 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2024 = T2025 || T1667;
  assign T2025 = T2026 || T1669;
  assign T2026 = T2027 || T1671;
  assign T2027 = T2028 || T1673;
  assign T2028 = T2029 || T1675;
  assign T2029 = T2030 || T1677;
  assign T2030 = T2031 || T1679;
  assign T2031 = T1682 || T1681;
  assign T2032 = T2118 | T2033;
  assign T2033 = State_1 & T2034;
  assign T2034 = {4'h8/* 8*/{T882}};
  assign T2035 = T2036 || T1696;
  assign T2036 = T2037 || T1698;
  assign T2037 = T2038 || T1700;
  assign T2038 = T2039 || T1702;
  assign T2039 = T2040 || T1704;
  assign T2040 = T2041 || T1706;
  assign T2041 = T2042 || T1708;
  assign T2042 = T2043 || T1710;
  assign T2043 = T2044 || T1711;
  assign T2044 = T2046 || T2045;
  assign T2045 = T830 && T882;
  assign T2046 = T2047 || T983;
  assign T2047 = T2049 || T2048;
  assign T2048 = T997 && T882;
  assign T2049 = T2050 || T1055;
  assign T2050 = T2052 || T2051;
  assign T2051 = T1069 && T882;
  assign T2052 = T2053 || T1127;
  assign T2053 = T2055 || T2054;
  assign T2054 = T1141 && T882;
  assign T2055 = T2056 || T1199;
  assign T2056 = T2058 || T2057;
  assign T2057 = T1213 && T882;
  assign T2058 = T2059 || T1271;
  assign T2059 = T2061 || T2060;
  assign T2060 = T1285 && T882;
  assign T2061 = T2062 || T1343;
  assign T2062 = T2064 || T2063;
  assign T2063 = T1357 && T882;
  assign T2064 = T2065 || T1415;
  assign T2065 = T2067 || T2066;
  assign T2066 = T1429 && T882;
  assign T2067 = T2068 || T1487;
  assign T2068 = T2070 || T2069;
  assign T2069 = T1501 && T882;
  assign T2070 = T883 || T2071;
  assign T2071 = T1504 && T128;
  assign T2072 = T2110 ? 8'hff/* 255*/ : T2073;
  assign T2073 = T2045 ? T2109 : T2074;
  assign T2074 = T983 ? T2108 : T2075;
  assign T2075 = T2048 ? T2107 : T2076;
  assign T2076 = T1055 ? T2106 : T2077;
  assign T2077 = T2051 ? T2105 : T2078;
  assign T2078 = T1127 ? T2104 : T2079;
  assign T2079 = T2054 ? T2103 : T2080;
  assign T2080 = T1199 ? T2102 : T2081;
  assign T2081 = T2057 ? T2101 : T2082;
  assign T2082 = T1271 ? T2100 : T2083;
  assign T2083 = T2060 ? T2099 : T2084;
  assign T2084 = T1343 ? T2098 : T2085;
  assign T2085 = T2063 ? T2097 : T2086;
  assign T2086 = T1415 ? T2096 : T2087;
  assign T2087 = T2066 ? T2095 : T2088;
  assign T2088 = T1487 ? T2094 : T2089;
  assign T2089 = T2069 ? T2093 : T2090;
  assign T2090 = T2071 ? T1529 : T2091;
  assign T2091 = T883 ? T2092 : State_1;
  assign T2092 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2093 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2094 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2095 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2096 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2097 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2098 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2099 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2100 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2101 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2102 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2103 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2104 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2105 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2106 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2107 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2108 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2109 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2110 = T2111 || T1696;
  assign T2111 = T2112 || T1698;
  assign T2112 = T2113 || T1700;
  assign T2113 = T2114 || T1702;
  assign T2114 = T2115 || T1704;
  assign T2115 = T2116 || T1706;
  assign T2116 = T2117 || T1708;
  assign T2117 = T1711 || T1710;
  assign T2118 = State_0 & T2119;
  assign T2119 = {4'h8/* 8*/{T888}};
  assign T2120 = T2121 || T1724;
  assign T2121 = T2122 || T1726;
  assign T2122 = T2123 || T1728;
  assign T2123 = T2124 || T1730;
  assign T2124 = T2125 || T1732;
  assign T2125 = T2126 || T1734;
  assign T2126 = T2127 || T1736;
  assign T2127 = T2128 || T1738;
  assign T2128 = T2129 || T1739;
  assign T2129 = T2131 || T2130;
  assign T2130 = T830 && T888;
  assign T2131 = T2132 || T990;
  assign T2132 = T2134 || T2133;
  assign T2133 = T997 && T888;
  assign T2134 = T2135 || T1062;
  assign T2135 = T2137 || T2136;
  assign T2136 = T1069 && T888;
  assign T2137 = T2138 || T1134;
  assign T2138 = T2140 || T2139;
  assign T2139 = T1141 && T888;
  assign T2140 = T2141 || T1206;
  assign T2141 = T2143 || T2142;
  assign T2142 = T1213 && T888;
  assign T2143 = T2144 || T1278;
  assign T2144 = T2146 || T2145;
  assign T2145 = T1285 && T888;
  assign T2146 = T2147 || T1350;
  assign T2147 = T2149 || T2148;
  assign T2148 = T1357 && T888;
  assign T2149 = T2150 || T1422;
  assign T2150 = T2152 || T2151;
  assign T2151 = T1429 && T888;
  assign T2152 = T2153 || T1494;
  assign T2153 = T2155 || T2154;
  assign T2154 = T1501 && T888;
  assign T2155 = T889 || T2156;
  assign T2156 = T1504 && T138;
  assign T2157 = T2195 ? 8'hff/* 255*/ : T2158;
  assign T2158 = T2130 ? T2194 : T2159;
  assign T2159 = T990 ? T2193 : T2160;
  assign T2160 = T2133 ? T2192 : T2161;
  assign T2161 = T1062 ? T2191 : T2162;
  assign T2162 = T2136 ? T2190 : T2163;
  assign T2163 = T1134 ? T2189 : T2164;
  assign T2164 = T2139 ? T2188 : T2165;
  assign T2165 = T1206 ? T2187 : T2166;
  assign T2166 = T2142 ? T2186 : T2167;
  assign T2167 = T1278 ? T2185 : T2168;
  assign T2168 = T2145 ? T2184 : T2169;
  assign T2169 = T1350 ? T2183 : T2170;
  assign T2170 = T2148 ? T2182 : T2171;
  assign T2171 = T1422 ? T2181 : T2172;
  assign T2172 = T2151 ? T2180 : T2173;
  assign T2173 = T1494 ? T2179 : T2174;
  assign T2174 = T2154 ? T2178 : T2175;
  assign T2175 = T2156 ? T1529 : T2176;
  assign T2176 = T889 ? T2177 : State_0;
  assign T2177 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2178 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2179 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2180 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2181 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2182 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2183 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2184 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2185 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2186 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2187 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2188 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2189 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2190 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2191 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2192 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2193 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2194 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2195 = T2196 || T1724;
  assign T2196 = T2197 || T1726;
  assign T2197 = T2198 || T1728;
  assign T2198 = T2199 || T1730;
  assign T2199 = T2200 || T1732;
  assign T2200 = T2201 || T1734;
  assign T2201 = T2202 || T1736;
  assign T2202 = T1739 || T1738;
  assign T2203 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2204 = T2205 || T1562;
  assign T2205 = T2206 || T1564;
  assign T2206 = T2207 || T1566;
  assign T2207 = T2208 || T1568;
  assign T2208 = T2209 || T1570;
  assign T2209 = T2210 || T1572;
  assign T2210 = T2211 || T1574;
  assign T2211 = T2212 || T1575;
  assign T2212 = T2214 || T2213;
  assign T2213 = T830 && T764;
  assign T2214 = T2215 || T944;
  assign T2215 = T2217 || T2216;
  assign T2216 = T997 && T764;
  assign T2217 = T2218 || T1016;
  assign T2218 = T2220 || T2219;
  assign T2219 = T1069 && T764;
  assign T2220 = T2221 || T1088;
  assign T2221 = T2223 || T2222;
  assign T2222 = T1141 && T764;
  assign T2223 = T2224 || T1160;
  assign T2224 = T2226 || T2225;
  assign T2225 = T1213 && T764;
  assign T2226 = T2227 || T1232;
  assign T2227 = T2229 || T2228;
  assign T2228 = T1285 && T764;
  assign T2229 = T2230 || T1304;
  assign T2230 = T2232 || T2231;
  assign T2231 = T1357 && T764;
  assign T2232 = T2233 || T1376;
  assign T2233 = T2235 || T2234;
  assign T2234 = T1429 && T764;
  assign T2235 = T2236 || T1448;
  assign T2236 = T2238 || T2237;
  assign T2237 = T1501 && T764;
  assign T2238 = T849 || T2239;
  assign T2239 = T1504 && T73;
  assign T2240 = T2278 ? 8'hff/* 255*/ : T2241;
  assign T2241 = T2213 ? T2277 : T2242;
  assign T2242 = T944 ? T2276 : T2243;
  assign T2243 = T2216 ? T2275 : T2244;
  assign T2244 = T1016 ? T2274 : T2245;
  assign T2245 = T2219 ? T2273 : T2246;
  assign T2246 = T1088 ? T2272 : T2247;
  assign T2247 = T2222 ? T2271 : T2248;
  assign T2248 = T1160 ? T2270 : T2249;
  assign T2249 = T2225 ? T2269 : T2250;
  assign T2250 = T1232 ? T2268 : T2251;
  assign T2251 = T2228 ? T2267 : T2252;
  assign T2252 = T1304 ? T2266 : T2253;
  assign T2253 = T2231 ? T2265 : T2254;
  assign T2254 = T1376 ? T2264 : T2255;
  assign T2255 = T2234 ? T2263 : T2256;
  assign T2256 = T1448 ? T2262 : T2257;
  assign T2257 = T2237 ? T2261 : T2258;
  assign T2258 = T2239 ? T1529 : T2259;
  assign T2259 = T849 ? T2260 : State_6;
  assign T2260 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2261 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2262 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2263 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2264 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2265 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2266 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2267 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2268 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2269 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2270 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2271 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2272 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2273 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2274 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2275 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2276 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2277 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2278 = T2279 || T763;
  assign T2279 = T2280 || T1562;
  assign T2280 = T2281 || T1564;
  assign T2281 = T2282 || T1566;
  assign T2282 = T2283 || T1568;
  assign T2283 = T2284 || T1570;
  assign T2284 = T2285 || T1572;
  assign T2285 = T1575 || T1574;
  assign T2286 = T2288 && T2287;
  assign T2287 = State_6 != 8'h0/* 0*/;
  assign T2288 = AllOffloadsReady && T2289;
  assign T2289 = T2290 == rThreadEncoder_io_chosen;
  assign T2290 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T2291 = subStateTh_5 == 1'h0/* 0*/;
  assign T2292 = T2296 ? 1'h1/* 1*/ : T2293;
  assign T2293 = T2294 ? 1'h0/* 0*/ : subStateTh_5;
  assign T2294 = T2295 == vThreadEncoder_io_chosen;
  assign T2295 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T2296 = T2298 && T2297;
  assign T2297 = State_5 != 8'hff/* 255*/;
  assign T2298 = T2300 && T2299;
  assign T2299 = State_5 != 8'h0/* 0*/;
  assign T2300 = AllOffloadsReady && T2301;
  assign T2301 = T2302 == rThreadEncoder_io_chosen;
  assign T2302 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T2303 = subStateTh_4 == 1'h0/* 0*/;
  assign T2304 = T2308 ? 1'h1/* 1*/ : T2305;
  assign T2305 = T2306 ? 1'h0/* 0*/ : subStateTh_4;
  assign T2306 = T2307 == vThreadEncoder_io_chosen;
  assign T2307 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T2308 = T2310 && T2309;
  assign T2309 = State_4 != 8'hff/* 255*/;
  assign T2310 = T2312 && T2311;
  assign T2311 = State_4 != 8'h0/* 0*/;
  assign T2312 = AllOffloadsReady && T2313;
  assign T2313 = T2314 == rThreadEncoder_io_chosen;
  assign T2314 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T2315 = subStateTh_3 == 1'h0/* 0*/;
  assign T2316 = T2320 ? 1'h1/* 1*/ : T2317;
  assign T2317 = T2318 ? 1'h0/* 0*/ : subStateTh_3;
  assign T2318 = T2319 == vThreadEncoder_io_chosen;
  assign T2319 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T2320 = T2322 && T2321;
  assign T2321 = State_3 != 8'hff/* 255*/;
  assign T2322 = T2324 && T2323;
  assign T2323 = State_3 != 8'h0/* 0*/;
  assign T2324 = AllOffloadsReady && T2325;
  assign T2325 = T2326 == rThreadEncoder_io_chosen;
  assign T2326 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T2327 = subStateTh_2 == 1'h0/* 0*/;
  assign T2328 = T2332 ? 1'h1/* 1*/ : T2329;
  assign T2329 = T2330 ? 1'h0/* 0*/ : subStateTh_2;
  assign T2330 = T2331 == vThreadEncoder_io_chosen;
  assign T2331 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T2332 = T2334 && T2333;
  assign T2333 = State_2 != 8'hff/* 255*/;
  assign T2334 = T2336 && T2335;
  assign T2335 = State_2 != 8'h0/* 0*/;
  assign T2336 = AllOffloadsReady && T2337;
  assign T2337 = T2338 == rThreadEncoder_io_chosen;
  assign T2338 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T2339 = subStateTh_1 == 1'h0/* 0*/;
  assign T2340 = T2344 ? 1'h1/* 1*/ : T2341;
  assign T2341 = T2342 ? 1'h0/* 0*/ : subStateTh_1;
  assign T2342 = T2343 == vThreadEncoder_io_chosen;
  assign T2343 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T2344 = T2346 && T2345;
  assign T2345 = State_1 != 8'hff/* 255*/;
  assign T2346 = T2348 && T2347;
  assign T2347 = State_1 != 8'h0/* 0*/;
  assign T2348 = AllOffloadsReady && T2349;
  assign T2349 = T2350 == rThreadEncoder_io_chosen;
  assign T2350 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T2351 = subStateTh_0 == 1'h0/* 0*/;
  assign T2352 = T2356 ? 1'h1/* 1*/ : T2353;
  assign T2353 = T2354 ? 1'h0/* 0*/ : subStateTh_0;
  assign T2354 = T2355 == vThreadEncoder_io_chosen;
  assign T2355 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T2356 = T2358 && T2357;
  assign T2357 = State_0 != 8'hff/* 255*/;
  assign T2358 = T2360 && T2359;
  assign T2359 = State_0 != 8'h0/* 0*/;
  assign T2360 = AllOffloadsReady && T2361;
  assign T2361 = T2362 == rThreadEncoder_io_chosen;
  assign T2362 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T2363 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2364 = T2367 | T2365;
  assign T2365 = State_6 & T2366;
  assign T2366 = {4'h8/* 8*/{T73}};
  assign T2367 = T2370 | T2368;
  assign T2368 = State_5 & T2369;
  assign T2369 = {4'h8/* 8*/{T84}};
  assign T2370 = T2373 | T2371;
  assign T2371 = State_4 & T2372;
  assign T2372 = {4'h8/* 8*/{T95}};
  assign T2373 = T2376 | T2374;
  assign T2374 = State_3 & T2375;
  assign T2375 = {4'h8/* 8*/{T106}};
  assign T2376 = T2379 | T2377;
  assign T2377 = State_2 & T2378;
  assign T2378 = {4'h8/* 8*/{T117}};
  assign T2379 = T2382 | T2380;
  assign T2380 = State_1 & T2381;
  assign T2381 = {4'h8/* 8*/{T128}};
  assign T2382 = State_0 & T2383;
  assign T2383 = {4'h8/* 8*/{T138}};
  assign T2384 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2385 = T2467 && T2386;
  assign T2386 = ! T2387;
  assign T2387 = T2398 | T2388;
  assign T2388 = dramBank7_valid_received_7 & T22;
  assign T2389 = T2395 && T2390;
  assign T2390 = dramBank7_valid_received_7 || T2391;
  assign T2391 = dramBank7Port_rep_valid && T2392;
  assign T2392 = dramBank7Port_rep_tag == T2393;
  assign T2393 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank7Port_rep_tag = mainOff_dramBank7_rep_tag;
  assign mainOff_dramBank7_req_tag = dramBank7Port_req_tag;
  assign dramBank7Port_req_tag = T2394;
  assign T2394 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank7Port_rep_valid = mainOff_dramBank7_rep_valid;
  assign T2395 = ! T2396;
  assign T2396 = T2397 == 5'h7/* 7*/;
  assign T2397 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2398 = T2408 | T2399;
  assign T2399 = dramBank7_valid_received_6 & T73;
  assign T2400 = T2405 && T2401;
  assign T2401 = dramBank7_valid_received_6 || T2402;
  assign T2402 = dramBank7Port_rep_valid && T2403;
  assign T2403 = dramBank7Port_rep_tag == T2404;
  assign T2404 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2405 = ! T2406;
  assign T2406 = T2407 == 5'h6/* 6*/;
  assign T2407 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2408 = T2418 | T2409;
  assign T2409 = dramBank7_valid_received_5 & T84;
  assign T2410 = T2415 && T2411;
  assign T2411 = dramBank7_valid_received_5 || T2412;
  assign T2412 = dramBank7Port_rep_valid && T2413;
  assign T2413 = dramBank7Port_rep_tag == T2414;
  assign T2414 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2415 = ! T2416;
  assign T2416 = T2417 == 5'h5/* 5*/;
  assign T2417 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2418 = T2428 | T2419;
  assign T2419 = dramBank7_valid_received_4 & T95;
  assign T2420 = T2425 && T2421;
  assign T2421 = dramBank7_valid_received_4 || T2422;
  assign T2422 = dramBank7Port_rep_valid && T2423;
  assign T2423 = dramBank7Port_rep_tag == T2424;
  assign T2424 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2425 = ! T2426;
  assign T2426 = T2427 == 5'h4/* 4*/;
  assign T2427 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2428 = T2438 | T2429;
  assign T2429 = dramBank7_valid_received_3 & T106;
  assign T2430 = T2435 && T2431;
  assign T2431 = dramBank7_valid_received_3 || T2432;
  assign T2432 = dramBank7Port_rep_valid && T2433;
  assign T2433 = dramBank7Port_rep_tag == T2434;
  assign T2434 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2435 = ! T2436;
  assign T2436 = T2437 == 5'h3/* 3*/;
  assign T2437 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2438 = T2448 | T2439;
  assign T2439 = dramBank7_valid_received_2 & T117;
  assign T2440 = T2445 && T2441;
  assign T2441 = dramBank7_valid_received_2 || T2442;
  assign T2442 = dramBank7Port_rep_valid && T2443;
  assign T2443 = dramBank7Port_rep_tag == T2444;
  assign T2444 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T2445 = ! T2446;
  assign T2446 = T2447 == 5'h2/* 2*/;
  assign T2447 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2448 = T2458 | T2449;
  assign T2449 = dramBank7_valid_received_1 & T128;
  assign T2450 = T2455 && T2451;
  assign T2451 = dramBank7_valid_received_1 || T2452;
  assign T2452 = dramBank7Port_rep_valid && T2453;
  assign T2453 = dramBank7Port_rep_tag == T2454;
  assign T2454 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T2455 = ! T2456;
  assign T2456 = T2457 == 5'h1/* 1*/;
  assign T2457 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2458 = dramBank7_valid_received_0 & T138;
  assign T2459 = T2464 && T2460;
  assign T2460 = dramBank7_valid_received_0 || T2461;
  assign T2461 = dramBank7Port_rep_valid && T2462;
  assign T2462 = dramBank7Port_rep_tag == T2463;
  assign T2463 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T2464 = ! T2465;
  assign T2465 = T2466 == 5'h0/* 0*/;
  assign T2466 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2467 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2468 = 5'h7/* 7*/ == T2469;
  assign T2469 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2470 = ! T2471;
  assign T2471 = T2472 == 5'h7/* 7*/;
  assign T2472 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2473 = T2474 || dramBank7_valid_received_7;
  assign T2474 = dramBank7Port_rep_valid && T2475;
  assign T2475 = dramBank7Port_rep_tag == T2476;
  assign T2476 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2477 = T2492 && T2478;
  assign T2478 = T2488 || T2479;
  assign T2479 = ! dramBank6PortHadValidRequest_7;
  assign T2480 = T2485 && T2481;
  assign T2481 = dramBank6PortHadValidRequest_7 || T2482;
  assign T2482 = T2483 && dramBank6Port_req_valid;
  assign T2483 = 5'h7/* 7*/ == T2484;
  assign T2484 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2485 = ! T2486;
  assign T2486 = T2487 == 5'h7/* 7*/;
  assign T2487 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2488 = T2489 || dramBank6_valid_received_7;
  assign T2489 = dramBank6Port_rep_valid && T2490;
  assign T2490 = dramBank6Port_rep_tag == T2491;
  assign T2491 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2492 = T2507 && T2493;
  assign T2493 = T2503 || T2494;
  assign T2494 = ! dramBank5PortHadValidRequest_7;
  assign T2495 = T2500 && T2496;
  assign T2496 = dramBank5PortHadValidRequest_7 || T2497;
  assign T2497 = T2498 && dramBank5Port_req_valid;
  assign T2498 = 5'h7/* 7*/ == T2499;
  assign T2499 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2500 = ! T2501;
  assign T2501 = T2502 == 5'h7/* 7*/;
  assign T2502 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2503 = T2504 || dramBank5_valid_received_7;
  assign T2504 = dramBank5Port_rep_valid && T2505;
  assign T2505 = dramBank5Port_rep_tag == T2506;
  assign T2506 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2507 = T2522 && T2508;
  assign T2508 = T2518 || T2509;
  assign T2509 = ! dramBank4PortHadValidRequest_7;
  assign T2510 = T2515 && T2511;
  assign T2511 = dramBank4PortHadValidRequest_7 || T2512;
  assign T2512 = T2513 && dramBank4Port_req_valid;
  assign T2513 = 5'h7/* 7*/ == T2514;
  assign T2514 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2515 = ! T2516;
  assign T2516 = T2517 == 5'h7/* 7*/;
  assign T2517 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2518 = T2519 || dramBank4_valid_received_7;
  assign T2519 = dramBank4Port_rep_valid && T2520;
  assign T2520 = dramBank4Port_rep_tag == T2521;
  assign T2521 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2522 = T2537 && T2523;
  assign T2523 = T2533 || T2524;
  assign T2524 = ! dramBank3PortHadValidRequest_7;
  assign T2525 = T2530 && T2526;
  assign T2526 = dramBank3PortHadValidRequest_7 || T2527;
  assign T2527 = T2528 && dramBank3Port_req_valid;
  assign T2528 = 5'h7/* 7*/ == T2529;
  assign T2529 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2530 = ! T2531;
  assign T2531 = T2532 == 5'h7/* 7*/;
  assign T2532 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2533 = T2534 || dramBank3_valid_received_7;
  assign T2534 = dramBank3Port_rep_valid && T2535;
  assign T2535 = dramBank3Port_rep_tag == T2536;
  assign T2536 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2537 = T2552 && T2538;
  assign T2538 = T2548 || T2539;
  assign T2539 = ! dramBank2PortHadValidRequest_7;
  assign T2540 = T2545 && T2541;
  assign T2541 = dramBank2PortHadValidRequest_7 || T2542;
  assign T2542 = T2543 && dramBank2Port_req_valid;
  assign T2543 = 5'h7/* 7*/ == T2544;
  assign T2544 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2545 = ! T2546;
  assign T2546 = T2547 == 5'h7/* 7*/;
  assign T2547 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2548 = T2549 || dramBank2_valid_received_7;
  assign T2549 = dramBank2Port_rep_valid && T2550;
  assign T2550 = dramBank2Port_rep_tag == T2551;
  assign T2551 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2552 = T2567 && T2553;
  assign T2553 = T2563 || T2554;
  assign T2554 = ! dramBank1PortHadValidRequest_7;
  assign T2555 = T2560 && T2556;
  assign T2556 = dramBank1PortHadValidRequest_7 || T2557;
  assign T2557 = T2558 && dramBank1Port_req_valid;
  assign T2558 = 5'h7/* 7*/ == T2559;
  assign T2559 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2560 = ! T2561;
  assign T2561 = T2562 == 5'h7/* 7*/;
  assign T2562 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2563 = T2564 || dramBank1_valid_received_7;
  assign T2564 = dramBank1Port_rep_valid && T2565;
  assign T2565 = dramBank1Port_rep_tag == T2566;
  assign T2566 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2567 = T2577 || T2568;
  assign T2568 = ! dramBank0PortHadValidRequest_7;
  assign T2569 = T2574 && T2570;
  assign T2570 = dramBank0PortHadValidRequest_7 || T2571;
  assign T2571 = T2572 && dramBank0Port_req_valid;
  assign T2572 = 5'h7/* 7*/ == T2573;
  assign T2573 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2574 = ! T2575;
  assign T2575 = T2576 == 5'h7/* 7*/;
  assign T2576 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2577 = T2578 || dramBank0_valid_received_7;
  assign T2578 = dramBank0Port_rep_valid && T2579;
  assign T2579 = dramBank0Port_rep_tag == T2580;
  assign T2580 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2581 = subStateTh_7 == 1'h1/* 1*/;
  assign T2582 = T2702 && AllOffloadsValid_6;
  assign AllOffloadsValid_6 = T2583;
  assign T2583 = T2598 && T2584;
  assign T2584 = T2594 || T2585;
  assign T2585 = ! dramBank7PortHadValidRequest_6;
  assign T2586 = T2591 && T2587;
  assign T2587 = dramBank7PortHadValidRequest_6 || T2588;
  assign T2588 = T2589 && dramBank7Port_req_valid;
  assign T2589 = 5'h6/* 6*/ == T2590;
  assign T2590 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2591 = ! T2592;
  assign T2592 = T2593 == 5'h6/* 6*/;
  assign T2593 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2594 = T2595 || dramBank7_valid_received_6;
  assign T2595 = dramBank7Port_rep_valid && T2596;
  assign T2596 = dramBank7Port_rep_tag == T2597;
  assign T2597 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2598 = T2613 && T2599;
  assign T2599 = T2609 || T2600;
  assign T2600 = ! dramBank6PortHadValidRequest_6;
  assign T2601 = T2606 && T2602;
  assign T2602 = dramBank6PortHadValidRequest_6 || T2603;
  assign T2603 = T2604 && dramBank6Port_req_valid;
  assign T2604 = 5'h6/* 6*/ == T2605;
  assign T2605 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2606 = ! T2607;
  assign T2607 = T2608 == 5'h6/* 6*/;
  assign T2608 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2609 = T2610 || dramBank6_valid_received_6;
  assign T2610 = dramBank6Port_rep_valid && T2611;
  assign T2611 = dramBank6Port_rep_tag == T2612;
  assign T2612 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2613 = T2628 && T2614;
  assign T2614 = T2624 || T2615;
  assign T2615 = ! dramBank5PortHadValidRequest_6;
  assign T2616 = T2621 && T2617;
  assign T2617 = dramBank5PortHadValidRequest_6 || T2618;
  assign T2618 = T2619 && dramBank5Port_req_valid;
  assign T2619 = 5'h6/* 6*/ == T2620;
  assign T2620 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2621 = ! T2622;
  assign T2622 = T2623 == 5'h6/* 6*/;
  assign T2623 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2624 = T2625 || dramBank5_valid_received_6;
  assign T2625 = dramBank5Port_rep_valid && T2626;
  assign T2626 = dramBank5Port_rep_tag == T2627;
  assign T2627 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2628 = T2643 && T2629;
  assign T2629 = T2639 || T2630;
  assign T2630 = ! dramBank4PortHadValidRequest_6;
  assign T2631 = T2636 && T2632;
  assign T2632 = dramBank4PortHadValidRequest_6 || T2633;
  assign T2633 = T2634 && dramBank4Port_req_valid;
  assign T2634 = 5'h6/* 6*/ == T2635;
  assign T2635 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2636 = ! T2637;
  assign T2637 = T2638 == 5'h6/* 6*/;
  assign T2638 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2639 = T2640 || dramBank4_valid_received_6;
  assign T2640 = dramBank4Port_rep_valid && T2641;
  assign T2641 = dramBank4Port_rep_tag == T2642;
  assign T2642 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2643 = T2658 && T2644;
  assign T2644 = T2654 || T2645;
  assign T2645 = ! dramBank3PortHadValidRequest_6;
  assign T2646 = T2651 && T2647;
  assign T2647 = dramBank3PortHadValidRequest_6 || T2648;
  assign T2648 = T2649 && dramBank3Port_req_valid;
  assign T2649 = 5'h6/* 6*/ == T2650;
  assign T2650 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2651 = ! T2652;
  assign T2652 = T2653 == 5'h6/* 6*/;
  assign T2653 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2654 = T2655 || dramBank3_valid_received_6;
  assign T2655 = dramBank3Port_rep_valid && T2656;
  assign T2656 = dramBank3Port_rep_tag == T2657;
  assign T2657 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2658 = T2673 && T2659;
  assign T2659 = T2669 || T2660;
  assign T2660 = ! dramBank2PortHadValidRequest_6;
  assign T2661 = T2666 && T2662;
  assign T2662 = dramBank2PortHadValidRequest_6 || T2663;
  assign T2663 = T2664 && dramBank2Port_req_valid;
  assign T2664 = 5'h6/* 6*/ == T2665;
  assign T2665 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2666 = ! T2667;
  assign T2667 = T2668 == 5'h6/* 6*/;
  assign T2668 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2669 = T2670 || dramBank2_valid_received_6;
  assign T2670 = dramBank2Port_rep_valid && T2671;
  assign T2671 = dramBank2Port_rep_tag == T2672;
  assign T2672 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2673 = T2688 && T2674;
  assign T2674 = T2684 || T2675;
  assign T2675 = ! dramBank1PortHadValidRequest_6;
  assign T2676 = T2681 && T2677;
  assign T2677 = dramBank1PortHadValidRequest_6 || T2678;
  assign T2678 = T2679 && dramBank1Port_req_valid;
  assign T2679 = 5'h6/* 6*/ == T2680;
  assign T2680 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2681 = ! T2682;
  assign T2682 = T2683 == 5'h6/* 6*/;
  assign T2683 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2684 = T2685 || dramBank1_valid_received_6;
  assign T2685 = dramBank1Port_rep_valid && T2686;
  assign T2686 = dramBank1Port_rep_tag == T2687;
  assign T2687 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2688 = T2698 || T2689;
  assign T2689 = ! dramBank0PortHadValidRequest_6;
  assign T2690 = T2695 && T2691;
  assign T2691 = dramBank0PortHadValidRequest_6 || T2692;
  assign T2692 = T2693 && dramBank0Port_req_valid;
  assign T2693 = 5'h6/* 6*/ == T2694;
  assign T2694 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2695 = ! T2696;
  assign T2696 = T2697 == 5'h6/* 6*/;
  assign T2697 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2698 = T2699 || dramBank0_valid_received_6;
  assign T2699 = dramBank0Port_rep_valid && T2700;
  assign T2700 = dramBank0Port_rep_tag == T2701;
  assign T2701 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2702 = subStateTh_6 == 1'h1/* 1*/;
  assign T2703 = T2823 && AllOffloadsValid_5;
  assign AllOffloadsValid_5 = T2704;
  assign T2704 = T2719 && T2705;
  assign T2705 = T2715 || T2706;
  assign T2706 = ! dramBank7PortHadValidRequest_5;
  assign T2707 = T2712 && T2708;
  assign T2708 = dramBank7PortHadValidRequest_5 || T2709;
  assign T2709 = T2710 && dramBank7Port_req_valid;
  assign T2710 = 5'h5/* 5*/ == T2711;
  assign T2711 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2712 = ! T2713;
  assign T2713 = T2714 == 5'h5/* 5*/;
  assign T2714 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2715 = T2716 || dramBank7_valid_received_5;
  assign T2716 = dramBank7Port_rep_valid && T2717;
  assign T2717 = dramBank7Port_rep_tag == T2718;
  assign T2718 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2719 = T2734 && T2720;
  assign T2720 = T2730 || T2721;
  assign T2721 = ! dramBank6PortHadValidRequest_5;
  assign T2722 = T2727 && T2723;
  assign T2723 = dramBank6PortHadValidRequest_5 || T2724;
  assign T2724 = T2725 && dramBank6Port_req_valid;
  assign T2725 = 5'h5/* 5*/ == T2726;
  assign T2726 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2727 = ! T2728;
  assign T2728 = T2729 == 5'h5/* 5*/;
  assign T2729 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2730 = T2731 || dramBank6_valid_received_5;
  assign T2731 = dramBank6Port_rep_valid && T2732;
  assign T2732 = dramBank6Port_rep_tag == T2733;
  assign T2733 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2734 = T2749 && T2735;
  assign T2735 = T2745 || T2736;
  assign T2736 = ! dramBank5PortHadValidRequest_5;
  assign T2737 = T2742 && T2738;
  assign T2738 = dramBank5PortHadValidRequest_5 || T2739;
  assign T2739 = T2740 && dramBank5Port_req_valid;
  assign T2740 = 5'h5/* 5*/ == T2741;
  assign T2741 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2742 = ! T2743;
  assign T2743 = T2744 == 5'h5/* 5*/;
  assign T2744 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2745 = T2746 || dramBank5_valid_received_5;
  assign T2746 = dramBank5Port_rep_valid && T2747;
  assign T2747 = dramBank5Port_rep_tag == T2748;
  assign T2748 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2749 = T2764 && T2750;
  assign T2750 = T2760 || T2751;
  assign T2751 = ! dramBank4PortHadValidRequest_5;
  assign T2752 = T2757 && T2753;
  assign T2753 = dramBank4PortHadValidRequest_5 || T2754;
  assign T2754 = T2755 && dramBank4Port_req_valid;
  assign T2755 = 5'h5/* 5*/ == T2756;
  assign T2756 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2757 = ! T2758;
  assign T2758 = T2759 == 5'h5/* 5*/;
  assign T2759 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2760 = T2761 || dramBank4_valid_received_5;
  assign T2761 = dramBank4Port_rep_valid && T2762;
  assign T2762 = dramBank4Port_rep_tag == T2763;
  assign T2763 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2764 = T2779 && T2765;
  assign T2765 = T2775 || T2766;
  assign T2766 = ! dramBank3PortHadValidRequest_5;
  assign T2767 = T2772 && T2768;
  assign T2768 = dramBank3PortHadValidRequest_5 || T2769;
  assign T2769 = T2770 && dramBank3Port_req_valid;
  assign T2770 = 5'h5/* 5*/ == T2771;
  assign T2771 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2772 = ! T2773;
  assign T2773 = T2774 == 5'h5/* 5*/;
  assign T2774 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2775 = T2776 || dramBank3_valid_received_5;
  assign T2776 = dramBank3Port_rep_valid && T2777;
  assign T2777 = dramBank3Port_rep_tag == T2778;
  assign T2778 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2779 = T2794 && T2780;
  assign T2780 = T2790 || T2781;
  assign T2781 = ! dramBank2PortHadValidRequest_5;
  assign T2782 = T2787 && T2783;
  assign T2783 = dramBank2PortHadValidRequest_5 || T2784;
  assign T2784 = T2785 && dramBank2Port_req_valid;
  assign T2785 = 5'h5/* 5*/ == T2786;
  assign T2786 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2787 = ! T2788;
  assign T2788 = T2789 == 5'h5/* 5*/;
  assign T2789 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2790 = T2791 || dramBank2_valid_received_5;
  assign T2791 = dramBank2Port_rep_valid && T2792;
  assign T2792 = dramBank2Port_rep_tag == T2793;
  assign T2793 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2794 = T2809 && T2795;
  assign T2795 = T2805 || T2796;
  assign T2796 = ! dramBank1PortHadValidRequest_5;
  assign T2797 = T2802 && T2798;
  assign T2798 = dramBank1PortHadValidRequest_5 || T2799;
  assign T2799 = T2800 && dramBank1Port_req_valid;
  assign T2800 = 5'h5/* 5*/ == T2801;
  assign T2801 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2802 = ! T2803;
  assign T2803 = T2804 == 5'h5/* 5*/;
  assign T2804 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2805 = T2806 || dramBank1_valid_received_5;
  assign T2806 = dramBank1Port_rep_valid && T2807;
  assign T2807 = dramBank1Port_rep_tag == T2808;
  assign T2808 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2809 = T2819 || T2810;
  assign T2810 = ! dramBank0PortHadValidRequest_5;
  assign T2811 = T2816 && T2812;
  assign T2812 = dramBank0PortHadValidRequest_5 || T2813;
  assign T2813 = T2814 && dramBank0Port_req_valid;
  assign T2814 = 5'h5/* 5*/ == T2815;
  assign T2815 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2816 = ! T2817;
  assign T2817 = T2818 == 5'h5/* 5*/;
  assign T2818 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2819 = T2820 || dramBank0_valid_received_5;
  assign T2820 = dramBank0Port_rep_valid && T2821;
  assign T2821 = dramBank0Port_rep_tag == T2822;
  assign T2822 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2823 = subStateTh_5 == 1'h1/* 1*/;
  assign T2824 = T2944 && AllOffloadsValid_4;
  assign AllOffloadsValid_4 = T2825;
  assign T2825 = T2840 && T2826;
  assign T2826 = T2836 || T2827;
  assign T2827 = ! dramBank7PortHadValidRequest_4;
  assign T2828 = T2833 && T2829;
  assign T2829 = dramBank7PortHadValidRequest_4 || T2830;
  assign T2830 = T2831 && dramBank7Port_req_valid;
  assign T2831 = 5'h4/* 4*/ == T2832;
  assign T2832 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2833 = ! T2834;
  assign T2834 = T2835 == 5'h4/* 4*/;
  assign T2835 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2836 = T2837 || dramBank7_valid_received_4;
  assign T2837 = dramBank7Port_rep_valid && T2838;
  assign T2838 = dramBank7Port_rep_tag == T2839;
  assign T2839 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2840 = T2855 && T2841;
  assign T2841 = T2851 || T2842;
  assign T2842 = ! dramBank6PortHadValidRequest_4;
  assign T2843 = T2848 && T2844;
  assign T2844 = dramBank6PortHadValidRequest_4 || T2845;
  assign T2845 = T2846 && dramBank6Port_req_valid;
  assign T2846 = 5'h4/* 4*/ == T2847;
  assign T2847 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2848 = ! T2849;
  assign T2849 = T2850 == 5'h4/* 4*/;
  assign T2850 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2851 = T2852 || dramBank6_valid_received_4;
  assign T2852 = dramBank6Port_rep_valid && T2853;
  assign T2853 = dramBank6Port_rep_tag == T2854;
  assign T2854 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2855 = T2870 && T2856;
  assign T2856 = T2866 || T2857;
  assign T2857 = ! dramBank5PortHadValidRequest_4;
  assign T2858 = T2863 && T2859;
  assign T2859 = dramBank5PortHadValidRequest_4 || T2860;
  assign T2860 = T2861 && dramBank5Port_req_valid;
  assign T2861 = 5'h4/* 4*/ == T2862;
  assign T2862 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2863 = ! T2864;
  assign T2864 = T2865 == 5'h4/* 4*/;
  assign T2865 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2866 = T2867 || dramBank5_valid_received_4;
  assign T2867 = dramBank5Port_rep_valid && T2868;
  assign T2868 = dramBank5Port_rep_tag == T2869;
  assign T2869 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2870 = T2885 && T2871;
  assign T2871 = T2881 || T2872;
  assign T2872 = ! dramBank4PortHadValidRequest_4;
  assign T2873 = T2878 && T2874;
  assign T2874 = dramBank4PortHadValidRequest_4 || T2875;
  assign T2875 = T2876 && dramBank4Port_req_valid;
  assign T2876 = 5'h4/* 4*/ == T2877;
  assign T2877 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2878 = ! T2879;
  assign T2879 = T2880 == 5'h4/* 4*/;
  assign T2880 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2881 = T2882 || dramBank4_valid_received_4;
  assign T2882 = dramBank4Port_rep_valid && T2883;
  assign T2883 = dramBank4Port_rep_tag == T2884;
  assign T2884 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2885 = T2900 && T2886;
  assign T2886 = T2896 || T2887;
  assign T2887 = ! dramBank3PortHadValidRequest_4;
  assign T2888 = T2893 && T2889;
  assign T2889 = dramBank3PortHadValidRequest_4 || T2890;
  assign T2890 = T2891 && dramBank3Port_req_valid;
  assign T2891 = 5'h4/* 4*/ == T2892;
  assign T2892 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2893 = ! T2894;
  assign T2894 = T2895 == 5'h4/* 4*/;
  assign T2895 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2896 = T2897 || dramBank3_valid_received_4;
  assign T2897 = dramBank3Port_rep_valid && T2898;
  assign T2898 = dramBank3Port_rep_tag == T2899;
  assign T2899 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2900 = T2915 && T2901;
  assign T2901 = T2911 || T2902;
  assign T2902 = ! dramBank2PortHadValidRequest_4;
  assign T2903 = T2908 && T2904;
  assign T2904 = dramBank2PortHadValidRequest_4 || T2905;
  assign T2905 = T2906 && dramBank2Port_req_valid;
  assign T2906 = 5'h4/* 4*/ == T2907;
  assign T2907 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2908 = ! T2909;
  assign T2909 = T2910 == 5'h4/* 4*/;
  assign T2910 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2911 = T2912 || dramBank2_valid_received_4;
  assign T2912 = dramBank2Port_rep_valid && T2913;
  assign T2913 = dramBank2Port_rep_tag == T2914;
  assign T2914 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2915 = T2930 && T2916;
  assign T2916 = T2926 || T2917;
  assign T2917 = ! dramBank1PortHadValidRequest_4;
  assign T2918 = T2923 && T2919;
  assign T2919 = dramBank1PortHadValidRequest_4 || T2920;
  assign T2920 = T2921 && dramBank1Port_req_valid;
  assign T2921 = 5'h4/* 4*/ == T2922;
  assign T2922 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2923 = ! T2924;
  assign T2924 = T2925 == 5'h4/* 4*/;
  assign T2925 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2926 = T2927 || dramBank1_valid_received_4;
  assign T2927 = dramBank1Port_rep_valid && T2928;
  assign T2928 = dramBank1Port_rep_tag == T2929;
  assign T2929 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2930 = T2940 || T2931;
  assign T2931 = ! dramBank0PortHadValidRequest_4;
  assign T2932 = T2937 && T2933;
  assign T2933 = dramBank0PortHadValidRequest_4 || T2934;
  assign T2934 = T2935 && dramBank0Port_req_valid;
  assign T2935 = 5'h4/* 4*/ == T2936;
  assign T2936 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2937 = ! T2938;
  assign T2938 = T2939 == 5'h4/* 4*/;
  assign T2939 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2940 = T2941 || dramBank0_valid_received_4;
  assign T2941 = dramBank0Port_rep_valid && T2942;
  assign T2942 = dramBank0Port_rep_tag == T2943;
  assign T2943 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2944 = subStateTh_4 == 1'h1/* 1*/;
  assign T2945 = T3065 && AllOffloadsValid_3;
  assign AllOffloadsValid_3 = T2946;
  assign T2946 = T2961 && T2947;
  assign T2947 = T2957 || T2948;
  assign T2948 = ! dramBank7PortHadValidRequest_3;
  assign T2949 = T2954 && T2950;
  assign T2950 = dramBank7PortHadValidRequest_3 || T2951;
  assign T2951 = T2952 && dramBank7Port_req_valid;
  assign T2952 = 5'h3/* 3*/ == T2953;
  assign T2953 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2954 = ! T2955;
  assign T2955 = T2956 == 5'h3/* 3*/;
  assign T2956 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2957 = T2958 || dramBank7_valid_received_3;
  assign T2958 = dramBank7Port_rep_valid && T2959;
  assign T2959 = dramBank7Port_rep_tag == T2960;
  assign T2960 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2961 = T2976 && T2962;
  assign T2962 = T2972 || T2963;
  assign T2963 = ! dramBank6PortHadValidRequest_3;
  assign T2964 = T2969 && T2965;
  assign T2965 = dramBank6PortHadValidRequest_3 || T2966;
  assign T2966 = T2967 && dramBank6Port_req_valid;
  assign T2967 = 5'h3/* 3*/ == T2968;
  assign T2968 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2969 = ! T2970;
  assign T2970 = T2971 == 5'h3/* 3*/;
  assign T2971 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2972 = T2973 || dramBank6_valid_received_3;
  assign T2973 = dramBank6Port_rep_valid && T2974;
  assign T2974 = dramBank6Port_rep_tag == T2975;
  assign T2975 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2976 = T2991 && T2977;
  assign T2977 = T2987 || T2978;
  assign T2978 = ! dramBank5PortHadValidRequest_3;
  assign T2979 = T2984 && T2980;
  assign T2980 = dramBank5PortHadValidRequest_3 || T2981;
  assign T2981 = T2982 && dramBank5Port_req_valid;
  assign T2982 = 5'h3/* 3*/ == T2983;
  assign T2983 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2984 = ! T2985;
  assign T2985 = T2986 == 5'h3/* 3*/;
  assign T2986 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2987 = T2988 || dramBank5_valid_received_3;
  assign T2988 = dramBank5Port_rep_valid && T2989;
  assign T2989 = dramBank5Port_rep_tag == T2990;
  assign T2990 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2991 = T3006 && T2992;
  assign T2992 = T3002 || T2993;
  assign T2993 = ! dramBank4PortHadValidRequest_3;
  assign T2994 = T2999 && T2995;
  assign T2995 = dramBank4PortHadValidRequest_3 || T2996;
  assign T2996 = T2997 && dramBank4Port_req_valid;
  assign T2997 = 5'h3/* 3*/ == T2998;
  assign T2998 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2999 = ! T3000;
  assign T3000 = T3001 == 5'h3/* 3*/;
  assign T3001 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3002 = T3003 || dramBank4_valid_received_3;
  assign T3003 = dramBank4Port_rep_valid && T3004;
  assign T3004 = dramBank4Port_rep_tag == T3005;
  assign T3005 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3006 = T3021 && T3007;
  assign T3007 = T3017 || T3008;
  assign T3008 = ! dramBank3PortHadValidRequest_3;
  assign T3009 = T3014 && T3010;
  assign T3010 = dramBank3PortHadValidRequest_3 || T3011;
  assign T3011 = T3012 && dramBank3Port_req_valid;
  assign T3012 = 5'h3/* 3*/ == T3013;
  assign T3013 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3014 = ! T3015;
  assign T3015 = T3016 == 5'h3/* 3*/;
  assign T3016 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3017 = T3018 || dramBank3_valid_received_3;
  assign T3018 = dramBank3Port_rep_valid && T3019;
  assign T3019 = dramBank3Port_rep_tag == T3020;
  assign T3020 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3021 = T3036 && T3022;
  assign T3022 = T3032 || T3023;
  assign T3023 = ! dramBank2PortHadValidRequest_3;
  assign T3024 = T3029 && T3025;
  assign T3025 = dramBank2PortHadValidRequest_3 || T3026;
  assign T3026 = T3027 && dramBank2Port_req_valid;
  assign T3027 = 5'h3/* 3*/ == T3028;
  assign T3028 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3029 = ! T3030;
  assign T3030 = T3031 == 5'h3/* 3*/;
  assign T3031 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3032 = T3033 || dramBank2_valid_received_3;
  assign T3033 = dramBank2Port_rep_valid && T3034;
  assign T3034 = dramBank2Port_rep_tag == T3035;
  assign T3035 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3036 = T3051 && T3037;
  assign T3037 = T3047 || T3038;
  assign T3038 = ! dramBank1PortHadValidRequest_3;
  assign T3039 = T3044 && T3040;
  assign T3040 = dramBank1PortHadValidRequest_3 || T3041;
  assign T3041 = T3042 && dramBank1Port_req_valid;
  assign T3042 = 5'h3/* 3*/ == T3043;
  assign T3043 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3044 = ! T3045;
  assign T3045 = T3046 == 5'h3/* 3*/;
  assign T3046 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3047 = T3048 || dramBank1_valid_received_3;
  assign T3048 = dramBank1Port_rep_valid && T3049;
  assign T3049 = dramBank1Port_rep_tag == T3050;
  assign T3050 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3051 = T3061 || T3052;
  assign T3052 = ! dramBank0PortHadValidRequest_3;
  assign T3053 = T3058 && T3054;
  assign T3054 = dramBank0PortHadValidRequest_3 || T3055;
  assign T3055 = T3056 && dramBank0Port_req_valid;
  assign T3056 = 5'h3/* 3*/ == T3057;
  assign T3057 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3058 = ! T3059;
  assign T3059 = T3060 == 5'h3/* 3*/;
  assign T3060 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3061 = T3062 || dramBank0_valid_received_3;
  assign T3062 = dramBank0Port_rep_valid && T3063;
  assign T3063 = dramBank0Port_rep_tag == T3064;
  assign T3064 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3065 = subStateTh_3 == 1'h1/* 1*/;
  assign T3066 = T3186 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T3067;
  assign T3067 = T3082 && T3068;
  assign T3068 = T3078 || T3069;
  assign T3069 = ! dramBank7PortHadValidRequest_2;
  assign T3070 = T3075 && T3071;
  assign T3071 = dramBank7PortHadValidRequest_2 || T3072;
  assign T3072 = T3073 && dramBank7Port_req_valid;
  assign T3073 = 5'h2/* 2*/ == T3074;
  assign T3074 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3075 = ! T3076;
  assign T3076 = T3077 == 5'h2/* 2*/;
  assign T3077 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3078 = T3079 || dramBank7_valid_received_2;
  assign T3079 = dramBank7Port_rep_valid && T3080;
  assign T3080 = dramBank7Port_rep_tag == T3081;
  assign T3081 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3082 = T3097 && T3083;
  assign T3083 = T3093 || T3084;
  assign T3084 = ! dramBank6PortHadValidRequest_2;
  assign T3085 = T3090 && T3086;
  assign T3086 = dramBank6PortHadValidRequest_2 || T3087;
  assign T3087 = T3088 && dramBank6Port_req_valid;
  assign T3088 = 5'h2/* 2*/ == T3089;
  assign T3089 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3090 = ! T3091;
  assign T3091 = T3092 == 5'h2/* 2*/;
  assign T3092 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3093 = T3094 || dramBank6_valid_received_2;
  assign T3094 = dramBank6Port_rep_valid && T3095;
  assign T3095 = dramBank6Port_rep_tag == T3096;
  assign T3096 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3097 = T3112 && T3098;
  assign T3098 = T3108 || T3099;
  assign T3099 = ! dramBank5PortHadValidRequest_2;
  assign T3100 = T3105 && T3101;
  assign T3101 = dramBank5PortHadValidRequest_2 || T3102;
  assign T3102 = T3103 && dramBank5Port_req_valid;
  assign T3103 = 5'h2/* 2*/ == T3104;
  assign T3104 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3105 = ! T3106;
  assign T3106 = T3107 == 5'h2/* 2*/;
  assign T3107 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3108 = T3109 || dramBank5_valid_received_2;
  assign T3109 = dramBank5Port_rep_valid && T3110;
  assign T3110 = dramBank5Port_rep_tag == T3111;
  assign T3111 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3112 = T3127 && T3113;
  assign T3113 = T3123 || T3114;
  assign T3114 = ! dramBank4PortHadValidRequest_2;
  assign T3115 = T3120 && T3116;
  assign T3116 = dramBank4PortHadValidRequest_2 || T3117;
  assign T3117 = T3118 && dramBank4Port_req_valid;
  assign T3118 = 5'h2/* 2*/ == T3119;
  assign T3119 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3120 = ! T3121;
  assign T3121 = T3122 == 5'h2/* 2*/;
  assign T3122 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3123 = T3124 || dramBank4_valid_received_2;
  assign T3124 = dramBank4Port_rep_valid && T3125;
  assign T3125 = dramBank4Port_rep_tag == T3126;
  assign T3126 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3127 = T3142 && T3128;
  assign T3128 = T3138 || T3129;
  assign T3129 = ! dramBank3PortHadValidRequest_2;
  assign T3130 = T3135 && T3131;
  assign T3131 = dramBank3PortHadValidRequest_2 || T3132;
  assign T3132 = T3133 && dramBank3Port_req_valid;
  assign T3133 = 5'h2/* 2*/ == T3134;
  assign T3134 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3135 = ! T3136;
  assign T3136 = T3137 == 5'h2/* 2*/;
  assign T3137 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3138 = T3139 || dramBank3_valid_received_2;
  assign T3139 = dramBank3Port_rep_valid && T3140;
  assign T3140 = dramBank3Port_rep_tag == T3141;
  assign T3141 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3142 = T3157 && T3143;
  assign T3143 = T3153 || T3144;
  assign T3144 = ! dramBank2PortHadValidRequest_2;
  assign T3145 = T3150 && T3146;
  assign T3146 = dramBank2PortHadValidRequest_2 || T3147;
  assign T3147 = T3148 && dramBank2Port_req_valid;
  assign T3148 = 5'h2/* 2*/ == T3149;
  assign T3149 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3150 = ! T3151;
  assign T3151 = T3152 == 5'h2/* 2*/;
  assign T3152 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3153 = T3154 || dramBank2_valid_received_2;
  assign T3154 = dramBank2Port_rep_valid && T3155;
  assign T3155 = dramBank2Port_rep_tag == T3156;
  assign T3156 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3157 = T3172 && T3158;
  assign T3158 = T3168 || T3159;
  assign T3159 = ! dramBank1PortHadValidRequest_2;
  assign T3160 = T3165 && T3161;
  assign T3161 = dramBank1PortHadValidRequest_2 || T3162;
  assign T3162 = T3163 && dramBank1Port_req_valid;
  assign T3163 = 5'h2/* 2*/ == T3164;
  assign T3164 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3165 = ! T3166;
  assign T3166 = T3167 == 5'h2/* 2*/;
  assign T3167 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3168 = T3169 || dramBank1_valid_received_2;
  assign T3169 = dramBank1Port_rep_valid && T3170;
  assign T3170 = dramBank1Port_rep_tag == T3171;
  assign T3171 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3172 = T3182 || T3173;
  assign T3173 = ! dramBank0PortHadValidRequest_2;
  assign T3174 = T3179 && T3175;
  assign T3175 = dramBank0PortHadValidRequest_2 || T3176;
  assign T3176 = T3177 && dramBank0Port_req_valid;
  assign T3177 = 5'h2/* 2*/ == T3178;
  assign T3178 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3179 = ! T3180;
  assign T3180 = T3181 == 5'h2/* 2*/;
  assign T3181 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3182 = T3183 || dramBank0_valid_received_2;
  assign T3183 = dramBank0Port_rep_valid && T3184;
  assign T3184 = dramBank0Port_rep_tag == T3185;
  assign T3185 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3186 = subStateTh_2 == 1'h1/* 1*/;
  assign T3187 = T3307 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T3188;
  assign T3188 = T3203 && T3189;
  assign T3189 = T3199 || T3190;
  assign T3190 = ! dramBank7PortHadValidRequest_1;
  assign T3191 = T3196 && T3192;
  assign T3192 = dramBank7PortHadValidRequest_1 || T3193;
  assign T3193 = T3194 && dramBank7Port_req_valid;
  assign T3194 = 5'h1/* 1*/ == T3195;
  assign T3195 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3196 = ! T3197;
  assign T3197 = T3198 == 5'h1/* 1*/;
  assign T3198 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3199 = T3200 || dramBank7_valid_received_1;
  assign T3200 = dramBank7Port_rep_valid && T3201;
  assign T3201 = dramBank7Port_rep_tag == T3202;
  assign T3202 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3203 = T3218 && T3204;
  assign T3204 = T3214 || T3205;
  assign T3205 = ! dramBank6PortHadValidRequest_1;
  assign T3206 = T3211 && T3207;
  assign T3207 = dramBank6PortHadValidRequest_1 || T3208;
  assign T3208 = T3209 && dramBank6Port_req_valid;
  assign T3209 = 5'h1/* 1*/ == T3210;
  assign T3210 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3211 = ! T3212;
  assign T3212 = T3213 == 5'h1/* 1*/;
  assign T3213 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3214 = T3215 || dramBank6_valid_received_1;
  assign T3215 = dramBank6Port_rep_valid && T3216;
  assign T3216 = dramBank6Port_rep_tag == T3217;
  assign T3217 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3218 = T3233 && T3219;
  assign T3219 = T3229 || T3220;
  assign T3220 = ! dramBank5PortHadValidRequest_1;
  assign T3221 = T3226 && T3222;
  assign T3222 = dramBank5PortHadValidRequest_1 || T3223;
  assign T3223 = T3224 && dramBank5Port_req_valid;
  assign T3224 = 5'h1/* 1*/ == T3225;
  assign T3225 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3226 = ! T3227;
  assign T3227 = T3228 == 5'h1/* 1*/;
  assign T3228 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3229 = T3230 || dramBank5_valid_received_1;
  assign T3230 = dramBank5Port_rep_valid && T3231;
  assign T3231 = dramBank5Port_rep_tag == T3232;
  assign T3232 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3233 = T3248 && T3234;
  assign T3234 = T3244 || T3235;
  assign T3235 = ! dramBank4PortHadValidRequest_1;
  assign T3236 = T3241 && T3237;
  assign T3237 = dramBank4PortHadValidRequest_1 || T3238;
  assign T3238 = T3239 && dramBank4Port_req_valid;
  assign T3239 = 5'h1/* 1*/ == T3240;
  assign T3240 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3241 = ! T3242;
  assign T3242 = T3243 == 5'h1/* 1*/;
  assign T3243 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3244 = T3245 || dramBank4_valid_received_1;
  assign T3245 = dramBank4Port_rep_valid && T3246;
  assign T3246 = dramBank4Port_rep_tag == T3247;
  assign T3247 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3248 = T3263 && T3249;
  assign T3249 = T3259 || T3250;
  assign T3250 = ! dramBank3PortHadValidRequest_1;
  assign T3251 = T3256 && T3252;
  assign T3252 = dramBank3PortHadValidRequest_1 || T3253;
  assign T3253 = T3254 && dramBank3Port_req_valid;
  assign T3254 = 5'h1/* 1*/ == T3255;
  assign T3255 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3256 = ! T3257;
  assign T3257 = T3258 == 5'h1/* 1*/;
  assign T3258 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3259 = T3260 || dramBank3_valid_received_1;
  assign T3260 = dramBank3Port_rep_valid && T3261;
  assign T3261 = dramBank3Port_rep_tag == T3262;
  assign T3262 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3263 = T3278 && T3264;
  assign T3264 = T3274 || T3265;
  assign T3265 = ! dramBank2PortHadValidRequest_1;
  assign T3266 = T3271 && T3267;
  assign T3267 = dramBank2PortHadValidRequest_1 || T3268;
  assign T3268 = T3269 && dramBank2Port_req_valid;
  assign T3269 = 5'h1/* 1*/ == T3270;
  assign T3270 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3271 = ! T3272;
  assign T3272 = T3273 == 5'h1/* 1*/;
  assign T3273 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3274 = T3275 || dramBank2_valid_received_1;
  assign T3275 = dramBank2Port_rep_valid && T3276;
  assign T3276 = dramBank2Port_rep_tag == T3277;
  assign T3277 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3278 = T3293 && T3279;
  assign T3279 = T3289 || T3280;
  assign T3280 = ! dramBank1PortHadValidRequest_1;
  assign T3281 = T3286 && T3282;
  assign T3282 = dramBank1PortHadValidRequest_1 || T3283;
  assign T3283 = T3284 && dramBank1Port_req_valid;
  assign T3284 = 5'h1/* 1*/ == T3285;
  assign T3285 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3286 = ! T3287;
  assign T3287 = T3288 == 5'h1/* 1*/;
  assign T3288 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3289 = T3290 || dramBank1_valid_received_1;
  assign T3290 = dramBank1Port_rep_valid && T3291;
  assign T3291 = dramBank1Port_rep_tag == T3292;
  assign T3292 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3293 = T3303 || T3294;
  assign T3294 = ! dramBank0PortHadValidRequest_1;
  assign T3295 = T3300 && T3296;
  assign T3296 = dramBank0PortHadValidRequest_1 || T3297;
  assign T3297 = T3298 && dramBank0Port_req_valid;
  assign T3298 = 5'h1/* 1*/ == T3299;
  assign T3299 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3300 = ! T3301;
  assign T3301 = T3302 == 5'h1/* 1*/;
  assign T3302 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3303 = T3304 || dramBank0_valid_received_1;
  assign T3304 = dramBank0Port_rep_valid && T3305;
  assign T3305 = dramBank0Port_rep_tag == T3306;
  assign T3306 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3307 = subStateTh_1 == 1'h1/* 1*/;
  assign T3308 = T3428 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T3309;
  assign T3309 = T3324 && T3310;
  assign T3310 = T3320 || T3311;
  assign T3311 = ! dramBank7PortHadValidRequest_0;
  assign T3312 = T3317 && T3313;
  assign T3313 = dramBank7PortHadValidRequest_0 || T3314;
  assign T3314 = T3315 && dramBank7Port_req_valid;
  assign T3315 = 5'h0/* 0*/ == T3316;
  assign T3316 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3317 = ! T3318;
  assign T3318 = T3319 == 5'h0/* 0*/;
  assign T3319 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3320 = T3321 || dramBank7_valid_received_0;
  assign T3321 = dramBank7Port_rep_valid && T3322;
  assign T3322 = dramBank7Port_rep_tag == T3323;
  assign T3323 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3324 = T3339 && T3325;
  assign T3325 = T3335 || T3326;
  assign T3326 = ! dramBank6PortHadValidRequest_0;
  assign T3327 = T3332 && T3328;
  assign T3328 = dramBank6PortHadValidRequest_0 || T3329;
  assign T3329 = T3330 && dramBank6Port_req_valid;
  assign T3330 = 5'h0/* 0*/ == T3331;
  assign T3331 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3332 = ! T3333;
  assign T3333 = T3334 == 5'h0/* 0*/;
  assign T3334 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3335 = T3336 || dramBank6_valid_received_0;
  assign T3336 = dramBank6Port_rep_valid && T3337;
  assign T3337 = dramBank6Port_rep_tag == T3338;
  assign T3338 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3339 = T3354 && T3340;
  assign T3340 = T3350 || T3341;
  assign T3341 = ! dramBank5PortHadValidRequest_0;
  assign T3342 = T3347 && T3343;
  assign T3343 = dramBank5PortHadValidRequest_0 || T3344;
  assign T3344 = T3345 && dramBank5Port_req_valid;
  assign T3345 = 5'h0/* 0*/ == T3346;
  assign T3346 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3347 = ! T3348;
  assign T3348 = T3349 == 5'h0/* 0*/;
  assign T3349 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3350 = T3351 || dramBank5_valid_received_0;
  assign T3351 = dramBank5Port_rep_valid && T3352;
  assign T3352 = dramBank5Port_rep_tag == T3353;
  assign T3353 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3354 = T3369 && T3355;
  assign T3355 = T3365 || T3356;
  assign T3356 = ! dramBank4PortHadValidRequest_0;
  assign T3357 = T3362 && T3358;
  assign T3358 = dramBank4PortHadValidRequest_0 || T3359;
  assign T3359 = T3360 && dramBank4Port_req_valid;
  assign T3360 = 5'h0/* 0*/ == T3361;
  assign T3361 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3362 = ! T3363;
  assign T3363 = T3364 == 5'h0/* 0*/;
  assign T3364 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3365 = T3366 || dramBank4_valid_received_0;
  assign T3366 = dramBank4Port_rep_valid && T3367;
  assign T3367 = dramBank4Port_rep_tag == T3368;
  assign T3368 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3369 = T3384 && T3370;
  assign T3370 = T3380 || T3371;
  assign T3371 = ! dramBank3PortHadValidRequest_0;
  assign T3372 = T3377 && T3373;
  assign T3373 = dramBank3PortHadValidRequest_0 || T3374;
  assign T3374 = T3375 && dramBank3Port_req_valid;
  assign T3375 = 5'h0/* 0*/ == T3376;
  assign T3376 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3377 = ! T3378;
  assign T3378 = T3379 == 5'h0/* 0*/;
  assign T3379 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3380 = T3381 || dramBank3_valid_received_0;
  assign T3381 = dramBank3Port_rep_valid && T3382;
  assign T3382 = dramBank3Port_rep_tag == T3383;
  assign T3383 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3384 = T3399 && T3385;
  assign T3385 = T3395 || T3386;
  assign T3386 = ! dramBank2PortHadValidRequest_0;
  assign T3387 = T3392 && T3388;
  assign T3388 = dramBank2PortHadValidRequest_0 || T3389;
  assign T3389 = T3390 && dramBank2Port_req_valid;
  assign T3390 = 5'h0/* 0*/ == T3391;
  assign T3391 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3392 = ! T3393;
  assign T3393 = T3394 == 5'h0/* 0*/;
  assign T3394 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3395 = T3396 || dramBank2_valid_received_0;
  assign T3396 = dramBank2Port_rep_valid && T3397;
  assign T3397 = dramBank2Port_rep_tag == T3398;
  assign T3398 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3399 = T3414 && T3400;
  assign T3400 = T3410 || T3401;
  assign T3401 = ! dramBank1PortHadValidRequest_0;
  assign T3402 = T3407 && T3403;
  assign T3403 = dramBank1PortHadValidRequest_0 || T3404;
  assign T3404 = T3405 && dramBank1Port_req_valid;
  assign T3405 = 5'h0/* 0*/ == T3406;
  assign T3406 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3407 = ! T3408;
  assign T3408 = T3409 == 5'h0/* 0*/;
  assign T3409 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3410 = T3411 || dramBank1_valid_received_0;
  assign T3411 = dramBank1Port_rep_valid && T3412;
  assign T3412 = dramBank1Port_rep_tag == T3413;
  assign T3413 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3414 = T3424 || T3415;
  assign T3415 = ! dramBank0PortHadValidRequest_0;
  assign T3416 = T3421 && T3417;
  assign T3417 = dramBank0PortHadValidRequest_0 || T3418;
  assign T3418 = T3419 && dramBank0Port_req_valid;
  assign T3419 = 5'h0/* 0*/ == T3420;
  assign T3420 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3421 = ! T3422;
  assign T3422 = T3423 == 5'h0/* 0*/;
  assign T3423 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3424 = T3425 || dramBank0_valid_received_0;
  assign T3425 = dramBank0Port_rep_valid && T3426;
  assign T3426 = dramBank0Port_rep_tag == T3427;
  assign T3427 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3428 = subStateTh_0 == 1'h1/* 1*/;
  assign T3429 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T3430 = T3431 || T1534;
  assign T3431 = T3432 || T1536;
  assign T3432 = T3433 || T1538;
  assign T3433 = T3434 || T1540;
  assign T3434 = T3435 || T1542;
  assign T3435 = T3436 || T1544;
  assign T3436 = T3437 || T1546;
  assign T3437 = T3438 || T1547;
  assign T3438 = T3440 || T3439;
  assign T3439 = T830 && T5;
  assign T3440 = T3441 || T936;
  assign T3441 = T3443 || T3442;
  assign T3442 = T997 && T5;
  assign T3443 = T3444 || T1008;
  assign T3444 = T3446 || T3445;
  assign T3445 = T1069 && T5;
  assign T3446 = T3447 || T1080;
  assign T3447 = T3449 || T3448;
  assign T3448 = T1141 && T5;
  assign T3449 = T3450 || T1152;
  assign T3450 = T3452 || T3451;
  assign T3451 = T1213 && T5;
  assign T3452 = T3453 || T1224;
  assign T3453 = T3455 || T3454;
  assign T3454 = T1285 && T5;
  assign T3455 = T3456 || T1296;
  assign T3456 = T3458 || T3457;
  assign T3457 = T1357 && T5;
  assign T3458 = T3459 || T1368;
  assign T3459 = T3461 || T3460;
  assign T3460 = T1429 && T5;
  assign T3461 = T3462 || T1440;
  assign T3462 = T3464 || T3463;
  assign T3463 = T1501 && T5;
  assign T3464 = T839 || T3465;
  assign T3465 = T1504 && T22;
  assign T3466 = T3504 ? 8'hff/* 255*/ : T3467;
  assign T3467 = T3439 ? T3503 : T3468;
  assign T3468 = T936 ? T3502 : T3469;
  assign T3469 = T3442 ? T3501 : T3470;
  assign T3470 = T1008 ? T3500 : T3471;
  assign T3471 = T3445 ? T3499 : T3472;
  assign T3472 = T1080 ? T3498 : T3473;
  assign T3473 = T3448 ? T3497 : T3474;
  assign T3474 = T1152 ? T3496 : T3475;
  assign T3475 = T3451 ? T3495 : T3476;
  assign T3476 = T1224 ? T3494 : T3477;
  assign T3477 = T3454 ? T3493 : T3478;
  assign T3478 = T1296 ? T3492 : T3479;
  assign T3479 = T3457 ? T3491 : T3480;
  assign T3480 = T1368 ? T3490 : T3481;
  assign T3481 = T3460 ? T3489 : T3482;
  assign T3482 = T1440 ? T3488 : T3483;
  assign T3483 = T3463 ? T3487 : T3484;
  assign T3484 = T3465 ? T1529 : T3485;
  assign T3485 = T839 ? T3486 : State_7;
  assign T3486 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T3487 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3488 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T3489 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3490 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T3491 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3492 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T3493 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T3495 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3496 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T3497 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3498 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T3499 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3500 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T3501 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3502 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T3503 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3504 = T3505 || T4;
  assign T3505 = T3506 || T1534;
  assign T3506 = T3507 || T1536;
  assign T3507 = T3508 || T1538;
  assign T3508 = T3509 || T1540;
  assign T3509 = T3510 || T1542;
  assign T3510 = T3511 || T1544;
  assign T3511 = T1547 || T1546;
  assign T3512 = subStateTh_7 == 1'h0/* 0*/;
  assign T3513 = T3515 && T3514;
  assign T3514 = State_6 == 8'h0/* 0*/;
  assign T3515 = subStateTh_6 == 1'h0/* 0*/;
  assign T3516 = T3518 && T3517;
  assign T3517 = State_5 == 8'h0/* 0*/;
  assign T3518 = subStateTh_5 == 1'h0/* 0*/;
  assign T3519 = T3521 && T3520;
  assign T3520 = State_4 == 8'h0/* 0*/;
  assign T3521 = subStateTh_4 == 1'h0/* 0*/;
  assign T3522 = T3524 && T3523;
  assign T3523 = State_3 == 8'h0/* 0*/;
  assign T3524 = subStateTh_3 == 1'h0/* 0*/;
  assign T3525 = T3527 && T3526;
  assign T3526 = State_2 == 8'h0/* 0*/;
  assign T3527 = subStateTh_2 == 1'h0/* 0*/;
  assign T3528 = T3530 && T3529;
  assign T3529 = State_1 == 8'h0/* 0*/;
  assign T3530 = subStateTh_1 == 1'h0/* 0*/;
  assign T3531 = T3533 && T3532;
  assign T3532 = State_0 == 8'h0/* 0*/;
  assign T3533 = subStateTh_0 == 1'h0/* 0*/;
  assign T3534 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign io_out_tag = T3535;
  assign T3535 = T3539 | T3536;
  assign T3536 = inputTag_7 & T3537;
  assign T3537 = {4'ha/* 10*/{T22}};
  assign T3538 = T839 ? io_in_tag : inputTag_7;
  assign T3539 = T3543 | T3540;
  assign T3540 = inputTag_6 & T3541;
  assign T3541 = {4'ha/* 10*/{T73}};
  assign T3542 = T849 ? io_in_tag : inputTag_6;
  assign T3543 = T3547 | T3544;
  assign T3544 = inputTag_5 & T3545;
  assign T3545 = {4'ha/* 10*/{T84}};
  assign T3546 = T855 ? io_in_tag : inputTag_5;
  assign T3547 = T3551 | T3548;
  assign T3548 = inputTag_4 & T3549;
  assign T3549 = {4'ha/* 10*/{T95}};
  assign T3550 = T862 ? io_in_tag : inputTag_4;
  assign T3551 = T3555 | T3552;
  assign T3552 = inputTag_3 & T3553;
  assign T3553 = {4'ha/* 10*/{T106}};
  assign T3554 = T869 ? io_in_tag : inputTag_3;
  assign T3555 = T3559 | T3556;
  assign T3556 = inputTag_2 & T3557;
  assign T3557 = {4'ha/* 10*/{T117}};
  assign T3558 = T876 ? io_in_tag : inputTag_2;
  assign T3559 = T3563 | T3560;
  assign T3560 = inputTag_1 & T3561;
  assign T3561 = {4'ha/* 10*/{T128}};
  assign T3562 = T883 ? io_in_tag : inputTag_1;
  assign T3563 = inputTag_0 & T3564;
  assign T3564 = {4'ha/* 10*/{T138}};
  assign T3565 = T889 ? io_in_tag : inputTag_0;
  assign io_out_valid = T3566;
  assign T3566 = T3568 && T3567;
  assign T3567 = T19 == 8'hff/* 255*/;
  assign T3568 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  RREncode_17 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T2351 ),
       .io_valid_1( T2339 ),
       .io_valid_2( T2327 ),
       .io_valid_3( T2315 ),
       .io_valid_4( T2303 ),
       .io_valid_5( T2291 ),
       .io_valid_6( T755 ),
       .io_valid_7( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T2363 ));
  RREncode_18 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T3308 ),
       .io_valid_1( T3187 ),
       .io_valid_2( T3066 ),
       .io_valid_3( T2945 ),
       .io_valid_4( T2824 ),
       .io_valid_5( T2703 ),
       .io_valid_6( T2582 ),
       .io_valid_7( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T3429 ));
  RREncode_19 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T3531 ),
       .io_valid_1( T3528 ),
       .io_valid_2( T3525 ),
       .io_valid_3( T3522 ),
       .io_valid_4( T3519 ),
       .io_valid_5( T3516 ),
       .io_valid_6( T3513 ),
       .io_valid_7( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T3534 ));

  always @(posedge clk) begin
    if(reset) begin
      State_7 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_7 <= T3466;
    end
    dramBank7PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_7 <= reset ? 1'h0/* 0*/ : T26;
    dramBank7PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T42;
    dramBank7_ready_received <= reset ? 1'h0/* 0*/ : T46;
    dramBank6_valid_received_7 <= reset ? 1'h0/* 0*/ : T62;
    dramBank6_valid_received_6 <= reset ? 1'h0/* 0*/ : T74;
    dramBank6_valid_received_5 <= reset ? 1'h0/* 0*/ : T85;
    dramBank6_valid_received_4 <= reset ? 1'h0/* 0*/ : T96;
    dramBank6_valid_received_3 <= reset ? 1'h0/* 0*/ : T107;
    dramBank6_valid_received_2 <= reset ? 1'h0/* 0*/ : T118;
    dramBank6_valid_received_1 <= reset ? 1'h0/* 0*/ : T129;
    dramBank6_valid_received_0 <= reset ? 1'h0/* 0*/ : T139;
    dramBank6PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T149;
    dramBank6_ready_received <= reset ? 1'h0/* 0*/ : T153;
    dramBank5_valid_received_7 <= reset ? 1'h0/* 0*/ : T169;
    dramBank5_valid_received_6 <= reset ? 1'h0/* 0*/ : T180;
    dramBank5_valid_received_5 <= reset ? 1'h0/* 0*/ : T190;
    dramBank5_valid_received_4 <= reset ? 1'h0/* 0*/ : T200;
    dramBank5_valid_received_3 <= reset ? 1'h0/* 0*/ : T210;
    dramBank5_valid_received_2 <= reset ? 1'h0/* 0*/ : T220;
    dramBank5_valid_received_1 <= reset ? 1'h0/* 0*/ : T230;
    dramBank5_valid_received_0 <= reset ? 1'h0/* 0*/ : T239;
    dramBank5PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T249;
    dramBank5_ready_received <= reset ? 1'h0/* 0*/ : T253;
    dramBank4_valid_received_7 <= reset ? 1'h0/* 0*/ : T269;
    dramBank4_valid_received_6 <= reset ? 1'h0/* 0*/ : T280;
    dramBank4_valid_received_5 <= reset ? 1'h0/* 0*/ : T290;
    dramBank4_valid_received_4 <= reset ? 1'h0/* 0*/ : T300;
    dramBank4_valid_received_3 <= reset ? 1'h0/* 0*/ : T310;
    dramBank4_valid_received_2 <= reset ? 1'h0/* 0*/ : T320;
    dramBank4_valid_received_1 <= reset ? 1'h0/* 0*/ : T330;
    dramBank4_valid_received_0 <= reset ? 1'h0/* 0*/ : T339;
    dramBank4PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T349;
    dramBank4_ready_received <= reset ? 1'h0/* 0*/ : T353;
    dramBank3_valid_received_7 <= reset ? 1'h0/* 0*/ : T369;
    dramBank3_valid_received_6 <= reset ? 1'h0/* 0*/ : T380;
    dramBank3_valid_received_5 <= reset ? 1'h0/* 0*/ : T390;
    dramBank3_valid_received_4 <= reset ? 1'h0/* 0*/ : T400;
    dramBank3_valid_received_3 <= reset ? 1'h0/* 0*/ : T410;
    dramBank3_valid_received_2 <= reset ? 1'h0/* 0*/ : T420;
    dramBank3_valid_received_1 <= reset ? 1'h0/* 0*/ : T430;
    dramBank3_valid_received_0 <= reset ? 1'h0/* 0*/ : T439;
    dramBank3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T449;
    dramBank3_ready_received <= reset ? 1'h0/* 0*/ : T453;
    dramBank2_valid_received_7 <= reset ? 1'h0/* 0*/ : T469;
    dramBank2_valid_received_6 <= reset ? 1'h0/* 0*/ : T480;
    dramBank2_valid_received_5 <= reset ? 1'h0/* 0*/ : T490;
    dramBank2_valid_received_4 <= reset ? 1'h0/* 0*/ : T500;
    dramBank2_valid_received_3 <= reset ? 1'h0/* 0*/ : T510;
    dramBank2_valid_received_2 <= reset ? 1'h0/* 0*/ : T520;
    dramBank2_valid_received_1 <= reset ? 1'h0/* 0*/ : T530;
    dramBank2_valid_received_0 <= reset ? 1'h0/* 0*/ : T539;
    dramBank2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T549;
    dramBank2_ready_received <= reset ? 1'h0/* 0*/ : T553;
    dramBank1_valid_received_7 <= reset ? 1'h0/* 0*/ : T569;
    dramBank1_valid_received_6 <= reset ? 1'h0/* 0*/ : T580;
    dramBank1_valid_received_5 <= reset ? 1'h0/* 0*/ : T590;
    dramBank1_valid_received_4 <= reset ? 1'h0/* 0*/ : T600;
    dramBank1_valid_received_3 <= reset ? 1'h0/* 0*/ : T610;
    dramBank1_valid_received_2 <= reset ? 1'h0/* 0*/ : T620;
    dramBank1_valid_received_1 <= reset ? 1'h0/* 0*/ : T630;
    dramBank1_valid_received_0 <= reset ? 1'h0/* 0*/ : T639;
    dramBank1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T649;
    dramBank1_ready_received <= reset ? 1'h0/* 0*/ : T653;
    dramBank0_valid_received_7 <= reset ? 1'h0/* 0*/ : T668;
    dramBank0_valid_received_6 <= reset ? 1'h0/* 0*/ : T679;
    dramBank0_valid_received_5 <= reset ? 1'h0/* 0*/ : T689;
    dramBank0_valid_received_4 <= reset ? 1'h0/* 0*/ : T699;
    dramBank0_valid_received_3 <= reset ? 1'h0/* 0*/ : T709;
    dramBank0_valid_received_2 <= reset ? 1'h0/* 0*/ : T719;
    dramBank0_valid_received_1 <= reset ? 1'h0/* 0*/ : T729;
    dramBank0_valid_received_0 <= reset ? 1'h0/* 0*/ : T738;
    dramBank0PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T748;
    dramBank0_ready_received <= reset ? 1'h0/* 0*/ : T752;
    subStateTh_6 <= reset ? 1'h0/* 0*/ : T756;
    if(reset) begin
      State_6 <= 8'h0/* 0*/;
    end else if(T762) begin
      State_6 <= T2240;
    end
    if(reset) begin
      State_5 <= 8'h0/* 0*/;
    end else if(T778) begin
      State_5 <= T1508;
    end
    if(T839) begin
      inputReg_7_addr <= T845;
    end
    if(T849) begin
      inputReg_6_addr <= T851;
    end
    if(T855) begin
      inputReg_5_addr <= T857;
    end
    if(T862) begin
      inputReg_4_addr <= T864;
    end
    if(T869) begin
      inputReg_3_addr <= T871;
    end
    if(T876) begin
      inputReg_2_addr <= T878;
    end
    if(T883) begin
      inputReg_1_addr <= T885;
    end
    if(T889) begin
      inputReg_0_addr <= T891;
    end
    if(reset) begin
      rb7RowAddr_7 <= 32'h0/* 0*/;
    end else if(T935) begin
      rb7RowAddr_7 <= T937;
    end
    if(reset) begin
      rb7RowAddr_6 <= 32'h0/* 0*/;
    end else if(T943) begin
      rb7RowAddr_6 <= T945;
    end
    if(reset) begin
      rb7RowAddr_5 <= 32'h0/* 0*/;
    end else if(T951) begin
      rb7RowAddr_5 <= T952;
    end
    if(reset) begin
      rb7RowAddr_4 <= 32'h0/* 0*/;
    end else if(T958) begin
      rb7RowAddr_4 <= T960;
    end
    if(reset) begin
      rb7RowAddr_3 <= 32'h0/* 0*/;
    end else if(T966) begin
      rb7RowAddr_3 <= T968;
    end
    if(reset) begin
      rb7RowAddr_2 <= 32'h0/* 0*/;
    end else if(T974) begin
      rb7RowAddr_2 <= T976;
    end
    if(reset) begin
      rb7RowAddr_1 <= 32'h0/* 0*/;
    end else if(T982) begin
      rb7RowAddr_1 <= T984;
    end
    if(reset) begin
      rb7RowAddr_0 <= 32'h0/* 0*/;
    end else if(T989) begin
      rb7RowAddr_0 <= T991;
    end
    if(reset) begin
      rb6RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1007) begin
      rb6RowAddr_7 <= T1009;
    end
    if(reset) begin
      rb6RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1015) begin
      rb6RowAddr_6 <= T1017;
    end
    if(reset) begin
      rb6RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1023) begin
      rb6RowAddr_5 <= T1024;
    end
    if(reset) begin
      rb6RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1030) begin
      rb6RowAddr_4 <= T1032;
    end
    if(reset) begin
      rb6RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1038) begin
      rb6RowAddr_3 <= T1040;
    end
    if(reset) begin
      rb6RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1046) begin
      rb6RowAddr_2 <= T1048;
    end
    if(reset) begin
      rb6RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1054) begin
      rb6RowAddr_1 <= T1056;
    end
    if(reset) begin
      rb6RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1061) begin
      rb6RowAddr_0 <= T1063;
    end
    if(reset) begin
      rb5RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1079) begin
      rb5RowAddr_7 <= T1081;
    end
    if(reset) begin
      rb5RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1087) begin
      rb5RowAddr_6 <= T1089;
    end
    if(reset) begin
      rb5RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1095) begin
      rb5RowAddr_5 <= T1096;
    end
    if(reset) begin
      rb5RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1102) begin
      rb5RowAddr_4 <= T1104;
    end
    if(reset) begin
      rb5RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1110) begin
      rb5RowAddr_3 <= T1112;
    end
    if(reset) begin
      rb5RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1118) begin
      rb5RowAddr_2 <= T1120;
    end
    if(reset) begin
      rb5RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1126) begin
      rb5RowAddr_1 <= T1128;
    end
    if(reset) begin
      rb5RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1133) begin
      rb5RowAddr_0 <= T1135;
    end
    if(reset) begin
      rb4RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1151) begin
      rb4RowAddr_7 <= T1153;
    end
    if(reset) begin
      rb4RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1159) begin
      rb4RowAddr_6 <= T1161;
    end
    if(reset) begin
      rb4RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1167) begin
      rb4RowAddr_5 <= T1168;
    end
    if(reset) begin
      rb4RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1174) begin
      rb4RowAddr_4 <= T1176;
    end
    if(reset) begin
      rb4RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1182) begin
      rb4RowAddr_3 <= T1184;
    end
    if(reset) begin
      rb4RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1190) begin
      rb4RowAddr_2 <= T1192;
    end
    if(reset) begin
      rb4RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1198) begin
      rb4RowAddr_1 <= T1200;
    end
    if(reset) begin
      rb4RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1205) begin
      rb4RowAddr_0 <= T1207;
    end
    if(reset) begin
      rb3RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1223) begin
      rb3RowAddr_7 <= T1225;
    end
    if(reset) begin
      rb3RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1231) begin
      rb3RowAddr_6 <= T1233;
    end
    if(reset) begin
      rb3RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1239) begin
      rb3RowAddr_5 <= T1240;
    end
    if(reset) begin
      rb3RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1246) begin
      rb3RowAddr_4 <= T1248;
    end
    if(reset) begin
      rb3RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1254) begin
      rb3RowAddr_3 <= T1256;
    end
    if(reset) begin
      rb3RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1262) begin
      rb3RowAddr_2 <= T1264;
    end
    if(reset) begin
      rb3RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1270) begin
      rb3RowAddr_1 <= T1272;
    end
    if(reset) begin
      rb3RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1277) begin
      rb3RowAddr_0 <= T1279;
    end
    if(reset) begin
      rb2RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1295) begin
      rb2RowAddr_7 <= T1297;
    end
    if(reset) begin
      rb2RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1303) begin
      rb2RowAddr_6 <= T1305;
    end
    if(reset) begin
      rb2RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1311) begin
      rb2RowAddr_5 <= T1312;
    end
    if(reset) begin
      rb2RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1318) begin
      rb2RowAddr_4 <= T1320;
    end
    if(reset) begin
      rb2RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1326) begin
      rb2RowAddr_3 <= T1328;
    end
    if(reset) begin
      rb2RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1334) begin
      rb2RowAddr_2 <= T1336;
    end
    if(reset) begin
      rb2RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1342) begin
      rb2RowAddr_1 <= T1344;
    end
    if(reset) begin
      rb2RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1349) begin
      rb2RowAddr_0 <= T1351;
    end
    if(reset) begin
      rb1RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1367) begin
      rb1RowAddr_7 <= T1369;
    end
    if(reset) begin
      rb1RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1375) begin
      rb1RowAddr_6 <= T1377;
    end
    if(reset) begin
      rb1RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1383) begin
      rb1RowAddr_5 <= T1384;
    end
    if(reset) begin
      rb1RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1390) begin
      rb1RowAddr_4 <= T1392;
    end
    if(reset) begin
      rb1RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1398) begin
      rb1RowAddr_3 <= T1400;
    end
    if(reset) begin
      rb1RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1406) begin
      rb1RowAddr_2 <= T1408;
    end
    if(reset) begin
      rb1RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1414) begin
      rb1RowAddr_1 <= T1416;
    end
    if(reset) begin
      rb1RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1421) begin
      rb1RowAddr_0 <= T1423;
    end
    if(reset) begin
      rb0RowAddr_7 <= 32'h1/* 1*/;
    end else if(T1439) begin
      rb0RowAddr_7 <= T1441;
    end
    if(reset) begin
      rb0RowAddr_6 <= 32'h1/* 1*/;
    end else if(T1447) begin
      rb0RowAddr_6 <= T1449;
    end
    if(reset) begin
      rb0RowAddr_5 <= 32'h1/* 1*/;
    end else if(T1455) begin
      rb0RowAddr_5 <= T1456;
    end
    if(reset) begin
      rb0RowAddr_4 <= 32'h1/* 1*/;
    end else if(T1462) begin
      rb0RowAddr_4 <= T1464;
    end
    if(reset) begin
      rb0RowAddr_3 <= 32'h1/* 1*/;
    end else if(T1470) begin
      rb0RowAddr_3 <= T1472;
    end
    if(reset) begin
      rb0RowAddr_2 <= 32'h1/* 1*/;
    end else if(T1478) begin
      rb0RowAddr_2 <= T1480;
    end
    if(reset) begin
      rb0RowAddr_1 <= 32'h1/* 1*/;
    end else if(T1486) begin
      rb0RowAddr_1 <= T1488;
    end
    if(reset) begin
      rb0RowAddr_0 <= 32'h1/* 1*/;
    end else if(T1493) begin
      rb0RowAddr_0 <= T1495;
    end
    if(reset) begin
      EmitReturnState_7 <= 8'h0/* 0*/;
    end else if(T1532) begin
      EmitReturnState_7 <= T1548;
    end
    if(reset) begin
      EmitReturnState_6 <= 8'h0/* 0*/;
    end else if(T1560) begin
      EmitReturnState_6 <= T1576;
    end
    if(reset) begin
      EmitReturnState_5 <= 8'h0/* 0*/;
    end else if(T1588) begin
      EmitReturnState_5 <= T1596;
    end
    if(reset) begin
      EmitReturnState_4 <= 8'h0/* 0*/;
    end else if(T1608) begin
      EmitReturnState_4 <= T1625;
    end
    if(reset) begin
      EmitReturnState_3 <= 8'h0/* 0*/;
    end else if(T1637) begin
      EmitReturnState_3 <= T1654;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T1666) begin
      EmitReturnState_2 <= T1683;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T1695) begin
      EmitReturnState_1 <= T1712;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T1723) begin
      EmitReturnState_0 <= T1740;
    end
    if(reset) begin
      State_4 <= 8'h0/* 0*/;
    end else if(T1777) begin
      State_4 <= T1814;
    end
    if(reset) begin
      State_3 <= 8'h0/* 0*/;
    end else if(T1863) begin
      State_3 <= T1900;
    end
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T1949) begin
      State_2 <= T1986;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T2035) begin
      State_1 <= T2072;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T2120) begin
      State_0 <= T2157;
    end
    subStateTh_5 <= reset ? 1'h0/* 0*/ : T2292;
    subStateTh_4 <= reset ? 1'h0/* 0*/ : T2304;
    subStateTh_3 <= reset ? 1'h0/* 0*/ : T2316;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T2328;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T2340;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T2352;
    dramBank7_valid_received_7 <= reset ? 1'h0/* 0*/ : T2389;
    dramBank7_valid_received_6 <= reset ? 1'h0/* 0*/ : T2400;
    dramBank7_valid_received_5 <= reset ? 1'h0/* 0*/ : T2410;
    dramBank7_valid_received_4 <= reset ? 1'h0/* 0*/ : T2420;
    dramBank7_valid_received_3 <= reset ? 1'h0/* 0*/ : T2430;
    dramBank7_valid_received_2 <= reset ? 1'h0/* 0*/ : T2440;
    dramBank7_valid_received_1 <= reset ? 1'h0/* 0*/ : T2450;
    dramBank7_valid_received_0 <= reset ? 1'h0/* 0*/ : T2459;
    dramBank6PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2480;
    dramBank5PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2495;
    dramBank4PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2510;
    dramBank3PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2525;
    dramBank2PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2540;
    dramBank1PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2555;
    dramBank0PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2569;
    dramBank7PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2586;
    dramBank6PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2601;
    dramBank5PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2616;
    dramBank4PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2631;
    dramBank3PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2646;
    dramBank2PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2661;
    dramBank1PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2676;
    dramBank0PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2690;
    dramBank7PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2707;
    dramBank6PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2722;
    dramBank5PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2737;
    dramBank4PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2752;
    dramBank3PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2767;
    dramBank2PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2782;
    dramBank1PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2797;
    dramBank0PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2811;
    dramBank7PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2828;
    dramBank6PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2843;
    dramBank5PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2858;
    dramBank4PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2873;
    dramBank3PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2888;
    dramBank2PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2903;
    dramBank1PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2918;
    dramBank0PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2932;
    dramBank7PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2949;
    dramBank6PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2964;
    dramBank5PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2979;
    dramBank4PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2994;
    dramBank3PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3009;
    dramBank2PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3024;
    dramBank1PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3039;
    dramBank0PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3053;
    dramBank7PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3070;
    dramBank6PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3085;
    dramBank5PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3100;
    dramBank4PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3115;
    dramBank3PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3130;
    dramBank2PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3145;
    dramBank1PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3160;
    dramBank0PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3174;
    dramBank7PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3191;
    dramBank6PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3206;
    dramBank5PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3221;
    dramBank4PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3236;
    dramBank3PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3251;
    dramBank2PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3266;
    dramBank1PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3281;
    dramBank0PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3295;
    dramBank7PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3312;
    dramBank6PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3327;
    dramBank5PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3342;
    dramBank4PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3357;
    dramBank3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3372;
    dramBank2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3387;
    dramBank1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3402;
    dramBank0PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3416;
    if(T839) begin
      inputTag_7 <= T3538;
    end
    if(T849) begin
      inputTag_6 <= T3542;
    end
    if(T855) begin
      inputTag_5 <= T3546;
    end
    if(T862) begin
      inputTag_4 <= T3550;
    end
    if(T869) begin
      inputTag_3 <= T3554;
    end
    if(T876) begin
      inputTag_2 <= T3558;
    end
    if(T883) begin
      inputTag_1 <= T3562;
    end
    if(T889) begin
      inputTag_0 <= T3565;
    end
  end
endmodule

module RREncode_20(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_21(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_22(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_20 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_21 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_22 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank1_req_ready,
    output mainOff_dramBank1_req_valid,
    output[31:0] mainOff_dramBank1_req_bits,
    output[9:0] mainOff_dramBank1_req_tag,
    output mainOff_dramBank1_rep_ready,
    input  mainOff_dramBank1_rep_valid,
    input [31:0] mainOff_dramBank1_rep_bits,
    input [9:0] mainOff_dramBank1_rep_tag,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire mainComp_mainOff_dramBank1_rep_ready;
  wire mainComp_mainOff_dramBank1_req_valid;
  wire[9:0] mainComp_mainOff_dramBank1_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank0_rep_ready;
  wire mainComp_mainOff_dramBank0_req_valid;
  wire[9:0] mainComp_mainOff_dramBank0_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank2_rep_ready = mainComp_mainOff_dramBank2_rep_ready;
  assign mainOff_dramBank2_req_valid = mainComp_mainOff_dramBank2_req_valid;
  assign mainOff_dramBank2_req_tag = mainComp_mainOff_dramBank2_req_tag;
  assign mainOff_dramBank1_rep_ready = mainComp_mainOff_dramBank1_rep_ready;
  assign mainOff_dramBank1_req_valid = mainComp_mainOff_dramBank1_req_valid;
  assign mainOff_dramBank1_req_tag = mainComp_mainOff_dramBank1_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  dram mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank0_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank0_req_valid( mainComp_mainOff_dramBank0_req_valid ),
       .mainOff_dramBank0_req_bits(  ),
       .mainOff_dramBank0_req_tag( mainComp_mainOff_dramBank0_req_tag ),
       .mainOff_dramBank0_rep_ready( mainComp_mainOff_dramBank0_rep_ready ),
       .mainOff_dramBank0_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank0_rep_bits(  ),
       .mainOff_dramBank0_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank1_req_ready( mainOff_dramBank1_req_ready ),
       .mainOff_dramBank1_req_valid( mainComp_mainOff_dramBank1_req_valid ),
       .mainOff_dramBank1_req_bits(  ),
       .mainOff_dramBank1_req_tag( mainComp_mainOff_dramBank1_req_tag ),
       .mainOff_dramBank1_rep_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .mainOff_dramBank1_rep_valid( mainOff_dramBank1_rep_valid ),
       .mainOff_dramBank1_rep_bits(  ),
       .mainOff_dramBank1_rep_tag( mainOff_dramBank1_rep_tag ),
       .mainOff_dramBank2_req_ready( mainOff_dramBank2_req_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( mainOff_dramBank2_rep_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( mainOff_dramBank2_rep_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank0_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank0_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank0_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_23(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_24(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_25(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_23 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_24 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_25 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank1_rep_ready;
  wire mainComp_mainOff_dramBank1_req_valid;
  wire[9:0] mainComp_mainOff_dramBank1_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank2_rep_ready = mainComp_mainOff_dramBank2_rep_ready;
  assign mainOff_dramBank2_req_valid = mainComp_mainOff_dramBank2_req_valid;
  assign mainOff_dramBank2_req_tag = mainComp_mainOff_dramBank2_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_7 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank1_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank1_req_valid( mainComp_mainOff_dramBank1_req_valid ),
       .mainOff_dramBank1_req_bits(  ),
       .mainOff_dramBank1_req_tag( mainComp_mainOff_dramBank1_req_tag ),
       .mainOff_dramBank1_rep_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .mainOff_dramBank1_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank1_rep_bits(  ),
       .mainOff_dramBank1_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank2_req_ready( mainOff_dramBank2_req_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( mainOff_dramBank2_rep_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( mainOff_dramBank2_rep_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank1_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank1_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_26(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_27(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_28(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_26 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_27 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_28 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_8 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank2_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_2 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank2_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank2_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_29(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_30(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_31(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_29 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_30 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_31 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_9 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank3_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_3 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank3_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank3_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_32(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_33(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_34(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_32 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_33 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_34 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_10 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank4_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank4_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank4_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_35(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_36(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_37(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_35 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_36 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_37 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_11 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank5_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_5 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank5_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank5_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_38(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_39(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_40(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_38 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_39 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_40 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_12 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank6_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_6 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank6_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank6_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_41(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_42(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_43(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire T0;
  wire sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_0;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  wire vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_0;
  wire T9;
  reg[0:0] subStateTh_0;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire rThreadEncoder_io_chosen;
  wire T19;
  wire AllOffloadsReady;
  wire T20;
  wire T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire[31:0] T31;
  reg[31:0] counter_0;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[7:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[7:0] T41;
  wire T42;
  wire[31:0] T43;
  wire[31:0] T44;
  wire[31:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire T75;
  wire[9:0] T76;
  wire[9:0] T77;
  reg[9:0] inputTag_0;
  wire[9:0] T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T1 = T75 && T2;
  assign T2 = State_0 == 8'h0/* 0*/;
  assign T3 = T26 || T4;
  assign T4 = T20 && T5;
  assign T5 = T6;
  assign T6 = T7[1'h0/* 0*/:1'h0/* 0*/];
  assign T7 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T9 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T9 = subStateTh_0 == 1'h1/* 1*/;
  assign T10 = T13 ? 1'h1/* 1*/ : T11;
  assign T11 = T12 ? 1'h0/* 0*/ : subStateTh_0;
  assign T12 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T13 = T15 && T14;
  assign T14 = State_0 != 8'hff/* 255*/;
  assign T15 = T17 && T16;
  assign T16 = State_0 != 8'h0/* 0*/;
  assign T17 = AllOffloadsReady && T18;
  assign T18 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign T19 = subStateTh_0 == 1'h0/* 0*/;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T20 = T25 && T21;
  assign T21 = T23 == T22;
  assign T22 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T23 = State_0 & T24;
  assign T24 = {4'h8/* 8*/{T5}};
  assign T25 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T26 = T46 || T27;
  assign T27 = T28 && T5;
  assign T28 = T34 && T29;
  assign T29 = T30 == 32'h0/* 0*/;
  assign T30 = counter_0 & T31;
  assign T31 = {6'h20/* 32*/{T5}};
  assign T32 = T38 || T33;
  assign T33 = T34 && T5;
  assign T34 = T37 && T35;
  assign T35 = T23 == T36;
  assign T36 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T37 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T38 = T39 && T5;
  assign T39 = T42 && T40;
  assign T40 = T23 == T41;
  assign T41 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T42 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T43 = T33 ? T45 : T44;
  assign T44 = T38 ? 32'ha/* 10*/ : counter_0;
  assign T45 = T30 - 32'h1/* 1*/;
  assign T46 = T47 || T38;
  assign T47 = T58 || T48;
  assign T48 = T52 && T49;
  assign T49 = T50;
  assign T50 = T51[1'h0/* 0*/:1'h0/* 0*/];
  assign T51 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T52 = T53 && io_out_ready;
  assign T53 = T57 && T54;
  assign T54 = T55 == 8'hff/* 255*/;
  assign T55 = State_0 & T56;
  assign T56 = {4'h8/* 8*/{T49}};
  assign T57 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T58 = T62 && T59;
  assign T59 = T60;
  assign T60 = T61[1'h0/* 0*/:1'h0/* 0*/];
  assign T61 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T62 = T63 && io_in_valid;
  assign T63 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T64 = T4 ? 8'hff/* 255*/ : T65;
  assign T65 = T27 ? T74 : T66;
  assign T66 = T38 ? T73 : T67;
  assign T67 = T48 ? T70 : T68;
  assign T68 = T58 ? T69 : State_0;
  assign T69 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T70 = EmitReturnState_0 & T71;
  assign T71 = {4'h8/* 8*/{T49}};
  assign T72 = T4 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T73 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T74 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign io_out_tag = T76;
  assign T76 = inputTag_0 & T77;
  assign T77 = {4'ha/* 10*/{T49}};
  assign T78 = T58 ? io_in_tag : inputTag_0;
  assign io_out_valid = T79;
  assign T79 = T81 && T80;
  assign T80 = T55 == 8'hff/* 255*/;
  assign T81 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_41 rThreadEncoder(
       .io_valid_0( T19 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_42 vThreadEncoder(
       .io_valid_0( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_43 sThreadEncoder(
       .io_valid_0( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_0 <= T64;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T10;
    if(T32) begin
      counter_0 <= T43;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_0 <= T72;
    end
    if(T58) begin
      inputTag_0 <= T78;
    end
  end
endmodule

module gOffloadedComponent_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire offComp_io_out_valid;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_13 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank7_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( offComp_io_out_tag ));
  dramBank_7 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank7_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank7_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_dram_req_valid;
  wire[31:0] mainComp_mainOff_dram_req_bits_addr;
  wire mainComp_io_out_valid;
  wire[127:0] mainComp_io_out_bits_data;
  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dram_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_dram_req_tag;
  wire offComp_io_out_valid;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_data = mainComp_io_out_bits_data;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_6 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data( mainComp_io_out_bits_data ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dram_req_ready( offComp_io_in_ready ),
       .mainOff_dram_req_valid( mainComp_mainOff_dram_req_valid ),
       .mainOff_dram_req_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .mainOff_dram_req_bits_rw(  ),
       .mainOff_dram_req_bits_cached(  ),
       .mainOff_dram_req_bits_data(  ),
       .mainOff_dram_req_bits_size(  ),
       .mainOff_dram_req_tag( mainComp_mainOff_dram_req_tag ),
       .mainOff_dram_rep_ready( mainComp_mainOff_dram_rep_ready ),
       .mainOff_dram_rep_valid( offComp_io_out_valid ),
       .mainOff_dram_rep_bits_data(  ),
       .mainOff_dram_rep_tag( offComp_io_out_tag ));
  gOffloadedComponent_14 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dram_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( mainComp_mainOff_dram_req_tag ),
       .io_out_ready( mainComp_mainOff_dram_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module prMemComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] generatedTop_io_out_tag;
  wire generatedTop_io_out_valid;
  wire[127:0] generatedTop_io_out_bits_data;
  wire generatedTop_io_in_ready;

  assign io_out_tag = generatedTop_io_out_tag;
  assign io_out_valid = generatedTop_io_out_valid;
  assign io_out_bits_data = generatedTop_io_out_bits_data;
  assign io_in_ready = generatedTop_io_in_ready;
  gOffloadedComponent_15 generatedTop(.clk(clk), .reset(reset),
       .io_in_ready( generatedTop_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( generatedTop_io_out_valid ),
       .io_out_bits_data( generatedTop_io_out_bits_data ),
       .io_out_tag( generatedTop_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_16(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire[9:0] offComp_io_out_tag;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire offComp_io_out_valid;
  wire[127:0] offComp_io_out_bits_data;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire mainComp_io_out_valid;
  wire mainComp_io_out_bits_done;
  wire[31:0] mainComp_io_out_bits_pageId;
  wire mainComp_mainOff_mem_req_valid;
  wire offComp_io_in_ready;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_done = mainComp_io_out_bits_done;
  assign io_out_bits_pageId = mainComp_io_out_bits_pageId;
  assign io_out_tag = mainComp_io_out_tag;
  gReplicatedComponent mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_done( mainComp_io_out_bits_done ),
       .io_out_bits_pageId( mainComp_io_out_bits_pageId ),
       .io_out_bits_rankUpdate(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( offComp_io_in_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( offComp_io_out_valid ),
       .mainOff_mem_rep_bits_data( offComp_io_out_bits_data ),
       .mainOff_mem_rep_tag( offComp_io_out_tag ));
  prMemComponent offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .io_in_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .io_in_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .io_in_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .io_in_tag( mainComp_mainOff_mem_req_tag ),
       .io_out_ready( mainComp_mainOff_mem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_data( offComp_io_out_bits_data ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_44(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_45(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_46(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateWriter(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_lock_req_ready,
    output mainOff_lock_req_valid,
    output[31:0] mainOff_lock_req_bits_id,
    output mainOff_lock_req_bits_op,
    output[9:0] mainOff_lock_req_tag,
    output mainOff_lock_rep_ready,
    input  mainOff_lock_rep_valid,
    input  mainOff_lock_rep_bits_out,
    input [9:0] mainOff_lock_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_1;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[4:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_1;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_1;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[4:0] T24;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_1;
  wire T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire AllOffloadsReady;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg[0:0] addPortHadReadyRequest;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg[0:0] add_ready_received;
  wire T46;
  wire T47;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire lockPort_req_valid;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[7:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  reg[0:0] lock_valid_received_1;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[9:0] T71;
  wire[9:0] lockPort_rep_tag;
  wire lockPort_rep_valid;
  wire T72;
  wire T73;
  wire[4:0] T74;
  wire T75;
  wire T76;
  reg[0:0] lock_valid_received_0;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[9:0] T81;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  reg[0:0] lockPortHadReadyRequest;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  reg[0:0] lock_ready_received;
  wire T91;
  wire T92;
  wire lockPort_req_ready;
  wire lockPort_rep_ready;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire memPort_req_valid;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire[7:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[7:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[7:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire[7:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mem_valid_received_1;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire[9:0] T125;
  wire[9:0] memPort_rep_tag;
  wire memPort_rep_valid;
  wire T126;
  wire T127;
  wire[4:0] T128;
  wire T129;
  reg[0:0] mem_valid_received_0;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[9:0] T134;
  wire T135;
  wire T136;
  wire[4:0] T137;
  wire T138;
  wire T139;
  reg[0:0] memPortHadReadyRequest;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg[0:0] mem_ready_received;
  wire T144;
  wire T145;
  wire memPort_req_ready;
  wire T146;
  wire T147;
  reg[0:0] subStateTh_0;
  wire T148;
  wire T149;
  wire T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  reg[7:0] State_0;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[7:0] T159;
  wire[7:0] T160;
  wire[7:0] T161;
  wire[7:0] T162;
  wire[7:0] T163;
  wire[7:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[7:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[7:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[7:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[7:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[7:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[7:0] T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  reg[0:0] inputReg_1_done;
  wire T214;
  wire T215;
  wire[1:0] T216;
  wire[4:0] T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  reg[0:0] inputReg_0_done;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire[7:0] T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[7:0] T241;
  wire[7:0] T242;
  wire[7:0] T243;
  wire[7:0] T244;
  wire[7:0] T245;
  wire[7:0] T246;
  wire[7:0] T247;
  wire[7:0] T248;
  wire[7:0] T249;
  wire[7:0] T250;
  wire[7:0] T251;
  wire[7:0] T252;
  wire[7:0] T253;
  wire[7:0] T254;
  wire[7:0] T255;
  reg[7:0] EmitReturnState_1;
  wire T256;
  wire T257;
  wire[7:0] T258;
  wire T259;
  wire[7:0] T260;
  wire[7:0] T261;
  reg[7:0] EmitReturnState_0;
  wire T262;
  wire[7:0] T263;
  wire T264;
  wire[7:0] T265;
  wire[7:0] T266;
  wire[7:0] T267;
  wire[7:0] T268;
  wire[7:0] T269;
  wire[7:0] T270;
  wire[7:0] T271;
  wire[7:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[1:0] T278;
  wire T279;
  wire[7:0] T280;
  wire[7:0] T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  reg[0:0] add_valid_received_1;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire[9:0] T291;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T292;
  wire addPort_rep_valid;
  wire T293;
  wire T294;
  wire[4:0] T295;
  wire T296;
  reg[0:0] add_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire T302;
  wire T303;
  wire[4:0] T304;
  wire T305;
  wire T306;
  wire[4:0] T307;
  wire T308;
  wire T309;
  wire[4:0] T310;
  wire T311;
  wire T312;
  wire T313;
  wire[9:0] T314;
  wire T315;
  wire T316;
  wire T317;
  reg[0:0] lockPortHadValidRequest_1;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire[4:0] T322;
  wire T323;
  wire T324;
  wire[4:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[9:0] T329;
  wire T330;
  wire T331;
  reg[0:0] memPortHadValidRequest_1;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire[4:0] T336;
  wire T337;
  wire T338;
  wire[4:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire[9:0] T343;
  wire T344;
  wire T345;
  wire AllOffloadsValid_0;
  wire T346;
  wire T347;
  wire T348;
  reg[0:0] addPortHadValidRequest_0;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[4:0] T353;
  wire T354;
  wire T355;
  wire[4:0] T356;
  wire T357;
  wire T358;
  wire T359;
  wire[9:0] T360;
  wire T361;
  wire T362;
  wire T363;
  reg[0:0] lockPortHadValidRequest_0;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[4:0] T368;
  wire T369;
  wire T370;
  wire[4:0] T371;
  wire T372;
  wire T373;
  wire T374;
  wire[9:0] T375;
  wire T376;
  wire T377;
  reg[0:0] memPortHadValidRequest_0;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[4:0] T382;
  wire T383;
  wire T384;
  wire[4:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire[9:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire[7:0] T411;
  wire[7:0] T412;
  wire[7:0] T413;
  wire[7:0] T414;
  wire[7:0] T415;
  wire[7:0] T416;
  wire[7:0] T417;
  wire[7:0] T418;
  wire[7:0] T419;
  wire[7:0] T420;
  wire[7:0] T421;
  wire[7:0] T422;
  wire[7:0] T423;
  wire[7:0] T424;
  wire[7:0] T425;
  wire[7:0] T426;
  wire[7:0] T427;
  wire[7:0] T428;
  wire[7:0] T429;
  wire[7:0] T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T437;
  wire[165:0] T438;
  wire[165:0] T439;
  wire[3:0] T440;
  wire[165:0] T441;
  wire[165:0] T442;
  wire[3:0] T443;
  wire[165:0] T444;
  wire[165:0] T445;
  wire[3:0] T446;
  wire[165:0] T447;
  wire[165:0] T448;
  wire[165:0] T449;
  wire[3:0] memReq4_size;
  wire[127:0] memReq4_data;
  wire[127:0] T450;
  wire[63:0] T451;
  wire[63:0] T452;
  wire[63:0] T453;
  reg[63:0] rank_1;
  wire T454;
  wire[127:0] T455;
  wire[127:0] T456;
  wire[127:0] T457;
  wire[127:0] T458;
  wire[127:0] T459;
  wire[127:0] T460;
  reg[127:0] memRep_1_data;
  wire T461;
  wire T462;
  wire T463;
  wire[127:0] T464;
  wire[127:0] T465;
  wire[127:0] memPortReplyValue;
  wire[127:0] T466;
  wire[127:0] T467;
  wire[127:0] T468;
  wire[127:0] T469;
  reg[127:0] memPortReplyStorage_1_data;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire[1024:0] T473;
  wire[127:0] T474;
  wire[127:0] memPort_rep_bits_data;
  wire[127:0] T475;
  wire[127:0] T476;
  reg[127:0] memPortReplyStorage_0_data;
  wire T477;
  wire T478;
  wire[127:0] T479;
  wire[127:0] T480;
  wire T481;
  wire T482;
  wire[9:0] T483;
  wire T484;
  wire T485;
  wire T486;
  wire[127:0] T487;
  wire[127:0] T488;
  reg[127:0] memRep_0_data;
  wire T489;
  wire T490;
  wire T491;
  wire[127:0] T492;
  wire T493;
  wire T494;
  wire T495;
  wire[127:0] T496;
  wire[63:0] addOut_out;
  wire[63:0] T497;
  wire[63:0] addPortReplyValue;
  wire[63:0] T498;
  wire[63:0] T499;
  wire[63:0] T500;
  wire[63:0] T501;
  reg[63:0] addPortReplyStorage_1_out;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire[1024:0] T505;
  wire[63:0] T506;
  wire[63:0] addPort_rep_bits_out;
  wire[63:0] T507;
  wire[63:0] T508;
  reg[63:0] addPortReplyStorage_0_out;
  wire T509;
  wire T510;
  wire[63:0] T511;
  wire[63:0] T512;
  wire T513;
  wire T514;
  wire[9:0] T515;
  wire[63:0] T516;
  wire[63:0] T517;
  reg[63:0] rank_0;
  wire T518;
  wire[127:0] T519;
  wire[127:0] T520;
  wire[127:0] T521;
  wire[127:0] T522;
  wire memReq4_cached;
  wire memReq4_rw;
  wire[31:0] memReq4_addr;
  wire[31:0] T523;
  wire[55:0] T524;
  wire[55:0] T525;
  wire[34:0] T526;
  wire[31:0] T527;
  wire[31:0] T528;
  wire[31:0] T529;
  reg[31:0] inputReg_1_pageId;
  wire[31:0] T530;
  wire[31:0] T531;
  wire[31:0] T532;
  reg[31:0] inputReg_0_pageId;
  wire[31:0] T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire T537;
  wire[127:0] T538;
  wire T539;
  wire T540;
  wire[31:0] T541;
  wire[165:0] T542;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T543;
  wire[55:0] T544;
  wire[55:0] T545;
  wire[34:0] T546;
  wire T547;
  wire T548;
  wire[7:0] T549;
  wire T550;
  wire[127:0] T551;
  wire T552;
  wire T553;
  wire[31:0] T554;
  wire[165:0] T555;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire[127:0] T556;
  wire[127:0] T557;
  wire[31:0] T558;
  wire[31:0] T559;
  wire[127:0] T560;
  wire[127:0] T561;
  wire[127:0] T562;
  wire[127:0] T563;
  wire[127:0] T564;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T565;
  wire[58:0] T566;
  wire[58:0] T567;
  wire[31:0] T568;
  wire T569;
  wire T570;
  wire[7:0] T571;
  wire T572;
  wire[127:0] T573;
  wire T574;
  wire T575;
  wire[31:0] T576;
  wire[165:0] T577;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T578;
  wire[58:0] T579;
  wire[58:0] T580;
  wire[31:0] T581;
  wire T582;
  wire T583;
  wire[7:0] T584;
  wire T585;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T586;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T587;
  wire memPort_req_bits_cached;
  wire T588;
  wire memPort_req_bits_rw;
  wire T589;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T590;
  wire[9:0] lockPort_req_tag;
  wire[9:0] T591;
  wire[9:0] T592;
  wire[9:0] T593;
  wire[9:0] T594;
  reg[9:0] inputTag_1;
  wire[9:0] T595;
  wire[9:0] T596;
  wire[9:0] T597;
  reg[9:0] inputTag_0;
  wire[9:0] T598;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T1 = T432 && T2;
  assign T2 = State_1 == 8'h0/* 0*/;
  assign T3 = T392 || T4;
  assign T4 = T157 && T5;
  assign T5 = T6[1'h1/* 1*/];
  assign T6 = T7[1'h1/* 1*/:1'h0/* 0*/];
  assign T7 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T344 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T9;
  assign T9 = T315 && T10;
  assign T10 = T311 || T11;
  assign T11 = ! addPortHadValidRequest_1;
  assign T12 = T308 && T13;
  assign T13 = addPortHadValidRequest_1 || T14;
  assign T14 = T306 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T283 && T16;
  assign T16 = T282 && T17;
  assign T17 = T19 == T18;
  assign T18 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T19 = T280 | T20;
  assign T20 = State_1 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23[1'h1/* 1*/];
  assign T23 = T24[1'h1/* 1*/:1'h0/* 0*/];
  assign T24 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_1 == 1'h0/* 0*/;
  assign T26 = T30 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_1;
  assign T28 = T29 == vThreadEncoder_io_chosen;
  assign T29 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T30 = T32 && T31;
  assign T31 = State_1 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_1 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = T36 == rThreadEncoder_io_chosen;
  assign T36 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign AllOffloadsReady = T37;
  assign T37 = T49 && T38;
  assign T38 = T45 || T39;
  assign T39 = T41 && T40;
  assign T40 = ! addPort_req_valid;
  assign T41 = ! addPortHadReadyRequest;
  assign T42 = T44 && T43;
  assign T43 = addPortHadReadyRequest || addPort_req_valid;
  assign T44 = ! AllOffloadsReady;
  assign T45 = addPort_req_ready || add_ready_received;
  assign T46 = T48 && T47;
  assign T47 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T48 = ! AllOffloadsReady;
  assign T49 = T94 && T50;
  assign T50 = T90 || T51;
  assign T51 = T86 && T52;
  assign T52 = ! lockPort_req_valid;
  assign lockPort_req_valid = T53;
  assign T53 = T63 && T54;
  assign T54 = T59 || T55;
  assign T55 = T58 && T56;
  assign T56 = T19 == T57;
  assign T57 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T58 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T59 = T62 && T60;
  assign T60 = T19 == T61;
  assign T61 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T63 = T85 && T64;
  assign T64 = ! T65;
  assign T65 = T75 | T66;
  assign T66 = lock_valid_received_1 & T22;
  assign T67 = T72 && T68;
  assign T68 = lock_valid_received_1 || T69;
  assign T69 = lockPort_rep_valid && T70;
  assign T70 = lockPort_rep_tag == T71;
  assign T71 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign lockPort_rep_tag = mainOff_lock_rep_tag;
  assign lockPort_rep_valid = mainOff_lock_rep_valid;
  assign T72 = ! T73;
  assign T73 = T74 == 5'h1/* 1*/;
  assign T74 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T75 = lock_valid_received_0 & T76;
  assign T76 = T23[1'h0/* 0*/];
  assign T77 = T82 && T78;
  assign T78 = lock_valid_received_0 || T79;
  assign T79 = lockPort_rep_valid && T80;
  assign T80 = lockPort_rep_tag == T81;
  assign T81 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T82 = ! T83;
  assign T83 = T84 == 5'h0/* 0*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T86 = ! lockPortHadReadyRequest;
  assign T87 = T89 && T88;
  assign T88 = lockPortHadReadyRequest || lockPort_req_valid;
  assign T89 = ! AllOffloadsReady;
  assign T90 = lockPort_req_ready || lock_ready_received;
  assign T91 = T93 && T92;
  assign T92 = lock_ready_received || lockPort_req_ready;
  assign lockPort_req_ready = mainOff_lock_req_ready;
  assign mainOff_lock_rep_ready = lockPort_rep_ready;
  assign lockPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_lock_req_valid = lockPort_req_valid;
  assign T93 = ! AllOffloadsReady;
  assign T94 = T143 || T95;
  assign T95 = T139 && T96;
  assign T96 = ! memPort_req_valid;
  assign memPort_req_valid = T97;
  assign T97 = T117 && T98;
  assign T98 = T103 || T99;
  assign T99 = T102 && T100;
  assign T100 = T19 == T101;
  assign T101 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T102 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T103 = T108 || T104;
  assign T104 = T107 && T105;
  assign T105 = T19 == T106;
  assign T106 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T107 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T108 = T113 || T109;
  assign T109 = T112 && T110;
  assign T110 = T19 == T111;
  assign T111 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T112 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T113 = T116 && T114;
  assign T114 = T19 == T115;
  assign T115 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T116 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T117 = T138 && T118;
  assign T118 = ! T119;
  assign T119 = T129 | T120;
  assign T120 = mem_valid_received_1 & T22;
  assign T121 = T126 && T122;
  assign T122 = mem_valid_received_1 || T123;
  assign T123 = memPort_rep_valid && T124;
  assign T124 = memPort_rep_tag == T125;
  assign T125 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T126 = ! T127;
  assign T127 = T128 == 5'h1/* 1*/;
  assign T128 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T129 = mem_valid_received_0 & T76;
  assign T130 = T135 && T131;
  assign T131 = mem_valid_received_0 || T132;
  assign T132 = memPort_rep_valid && T133;
  assign T133 = memPort_rep_tag == T134;
  assign T134 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T135 = ! T136;
  assign T136 = T137 == 5'h0/* 0*/;
  assign T137 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T138 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T139 = ! memPortHadReadyRequest;
  assign T140 = T142 && T141;
  assign T141 = memPortHadReadyRequest || memPort_req_valid;
  assign T142 = ! AllOffloadsReady;
  assign T143 = memPort_req_ready || mem_ready_received;
  assign T144 = T146 && T145;
  assign T145 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign mainOff_mem_req_valid = memPort_req_valid;
  assign T146 = ! AllOffloadsReady;
  assign T147 = subStateTh_0 == 1'h0/* 0*/;
  assign T148 = T152 ? 1'h1/* 1*/ : T149;
  assign T149 = T150 ? 1'h0/* 0*/ : subStateTh_0;
  assign T150 = T151 == vThreadEncoder_io_chosen;
  assign T151 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T152 = T274 && T153;
  assign T153 = State_0 != 8'hff/* 255*/;
  assign T154 = T166 || T155;
  assign T155 = T157 && T156;
  assign T156 = T6[1'h0/* 0*/];
  assign T157 = T165 && T158;
  assign T158 = T160 == T159;
  assign T159 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T160 = T163 | T161;
  assign T161 = State_1 & T162;
  assign T162 = {4'h8/* 8*/{T5}};
  assign T163 = State_0 & T164;
  assign T164 = {4'h8/* 8*/{T156}};
  assign T165 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T166 = T172 || T167;
  assign T167 = T168 && T156;
  assign T168 = T171 && T169;
  assign T169 = T160 == T170;
  assign T170 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T171 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T172 = T178 || T173;
  assign T173 = T174 && T156;
  assign T174 = T177 && T175;
  assign T175 = T160 == T176;
  assign T176 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T177 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T178 = T184 || T179;
  assign T179 = T180 && T156;
  assign T180 = T183 && T181;
  assign T181 = T160 == T182;
  assign T182 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T183 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T184 = T190 || T185;
  assign T185 = T186 && T156;
  assign T186 = T189 && T187;
  assign T187 = T160 == T188;
  assign T188 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T189 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T190 = T196 || T191;
  assign T191 = T192 && T156;
  assign T192 = T195 && T193;
  assign T193 = T160 == T194;
  assign T194 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T195 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T196 = T202 || T197;
  assign T197 = T198 && T156;
  assign T198 = T201 && T199;
  assign T199 = T160 == T200;
  assign T200 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T201 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T202 = T208 || T203;
  assign T203 = T204 && T156;
  assign T204 = T207 && T205;
  assign T205 = T160 == T206;
  assign T206 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T207 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T208 = T232 || T209;
  assign T209 = T210 && T156;
  assign T210 = T228 && T211;
  assign T211 = ! T212;
  assign T212 = T224 | T213;
  assign T213 = inputReg_1_done & T5;
  assign T214 = T218 && T215;
  assign T215 = T216[1'h1/* 1*/];
  assign T216 = T217[1'h1/* 1*/:1'h0/* 0*/];
  assign T217 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T218 = T222 && io_in_valid;
  assign io_out_valid = T219;
  assign T219 = T221 && T220;
  assign T220 = T19 == 8'hff/* 255*/;
  assign T221 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T222 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T223 = T214 ? io_in_bits_done : inputReg_1_done;
  assign T224 = inputReg_0_done & T156;
  assign T225 = T218 && T226;
  assign T226 = T216[1'h0/* 0*/];
  assign T227 = T225 ? io_in_bits_done : inputReg_0_done;
  assign T228 = T231 && T229;
  assign T229 = T160 == T230;
  assign T230 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T231 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T232 = T235 || T233;
  assign T233 = T234 && T156;
  assign T234 = T228 && T212;
  assign T235 = T225 || T236;
  assign T236 = T237 && T76;
  assign T237 = T238 && io_out_ready;
  assign T238 = T240 && T239;
  assign T239 = T19 == 8'hff/* 255*/;
  assign T240 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T241 = T273 ? 8'hff/* 255*/ : T242;
  assign T242 = T173 ? T272 : T243;
  assign T243 = T179 ? T271 : T244;
  assign T244 = T185 ? T270 : T245;
  assign T245 = T191 ? T269 : T246;
  assign T246 = T197 ? T268 : T247;
  assign T247 = T203 ? T267 : T248;
  assign T248 = T209 ? T266 : T249;
  assign T249 = T233 ? T265 : T250;
  assign T250 = T236 ? T253 : T251;
  assign T251 = T225 ? T252 : State_0;
  assign T252 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T253 = T260 | T254;
  assign T254 = EmitReturnState_1 & T255;
  assign T255 = {4'h8/* 8*/{T22}};
  assign T256 = T257 || T4;
  assign T257 = T168 && T5;
  assign T258 = T259 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T259 = T257 || T4;
  assign T260 = EmitReturnState_0 & T261;
  assign T261 = {4'h8/* 8*/{T76}};
  assign T262 = T167 || T155;
  assign T263 = T264 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T264 = T167 || T155;
  assign T265 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T266 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T267 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T268 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T269 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T270 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T271 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T272 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T273 = T167 || T155;
  assign T274 = T276 && T275;
  assign T275 = State_0 != 8'h0/* 0*/;
  assign T276 = AllOffloadsReady && T277;
  assign T277 = T278 == rThreadEncoder_io_chosen;
  assign T278 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T279 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T280 = State_0 & T281;
  assign T281 = {4'h8/* 8*/{T76}};
  assign T282 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T283 = T305 && T284;
  assign T284 = ! T285;
  assign T285 = T296 | T286;
  assign T286 = add_valid_received_1 & T22;
  assign T287 = T293 && T288;
  assign T288 = add_valid_received_1 || T289;
  assign T289 = addPort_rep_valid && T290;
  assign T290 = addPort_rep_tag == T291;
  assign T291 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T292;
  assign T292 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T293 = ! T294;
  assign T294 = T295 == 5'h1/* 1*/;
  assign T295 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T296 = add_valid_received_0 & T76;
  assign T297 = T302 && T298;
  assign T298 = add_valid_received_0 || T299;
  assign T299 = addPort_rep_valid && T300;
  assign T300 = addPort_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T302 = ! T303;
  assign T303 = T304 == 5'h0/* 0*/;
  assign T304 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T305 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T306 = 5'h1/* 1*/ == T307;
  assign T307 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T308 = ! T309;
  assign T309 = T310 == 5'h1/* 1*/;
  assign T310 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T311 = T312 || add_valid_received_1;
  assign T312 = addPort_rep_valid && T313;
  assign T313 = addPort_rep_tag == T314;
  assign T314 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T315 = T330 && T316;
  assign T316 = T326 || T317;
  assign T317 = ! lockPortHadValidRequest_1;
  assign T318 = T323 && T319;
  assign T319 = lockPortHadValidRequest_1 || T320;
  assign T320 = T321 && lockPort_req_valid;
  assign T321 = 5'h1/* 1*/ == T322;
  assign T322 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T323 = ! T324;
  assign T324 = T325 == 5'h1/* 1*/;
  assign T325 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T326 = T327 || lock_valid_received_1;
  assign T327 = lockPort_rep_valid && T328;
  assign T328 = lockPort_rep_tag == T329;
  assign T329 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T330 = T340 || T331;
  assign T331 = ! memPortHadValidRequest_1;
  assign T332 = T337 && T333;
  assign T333 = memPortHadValidRequest_1 || T334;
  assign T334 = T335 && memPort_req_valid;
  assign T335 = 5'h1/* 1*/ == T336;
  assign T336 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T337 = ! T338;
  assign T338 = T339 == 5'h1/* 1*/;
  assign T339 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T340 = T341 || mem_valid_received_1;
  assign T341 = memPort_rep_valid && T342;
  assign T342 = memPort_rep_tag == T343;
  assign T343 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T344 = subStateTh_1 == 1'h1/* 1*/;
  assign T345 = T390 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T346;
  assign T346 = T361 && T347;
  assign T347 = T357 || T348;
  assign T348 = ! addPortHadValidRequest_0;
  assign T349 = T354 && T350;
  assign T350 = addPortHadValidRequest_0 || T351;
  assign T351 = T352 && addPort_req_valid;
  assign T352 = 5'h0/* 0*/ == T353;
  assign T353 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T354 = ! T355;
  assign T355 = T356 == 5'h0/* 0*/;
  assign T356 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T357 = T358 || add_valid_received_0;
  assign T358 = addPort_rep_valid && T359;
  assign T359 = addPort_rep_tag == T360;
  assign T360 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T361 = T376 && T362;
  assign T362 = T372 || T363;
  assign T363 = ! lockPortHadValidRequest_0;
  assign T364 = T369 && T365;
  assign T365 = lockPortHadValidRequest_0 || T366;
  assign T366 = T367 && lockPort_req_valid;
  assign T367 = 5'h0/* 0*/ == T368;
  assign T368 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T369 = ! T370;
  assign T370 = T371 == 5'h0/* 0*/;
  assign T371 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T372 = T373 || lock_valid_received_0;
  assign T373 = lockPort_rep_valid && T374;
  assign T374 = lockPort_rep_tag == T375;
  assign T375 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T376 = T386 || T377;
  assign T377 = ! memPortHadValidRequest_0;
  assign T378 = T383 && T379;
  assign T379 = memPortHadValidRequest_0 || T380;
  assign T380 = T381 && memPort_req_valid;
  assign T381 = 5'h0/* 0*/ == T382;
  assign T382 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T383 = ! T384;
  assign T384 = T385 == 5'h0/* 0*/;
  assign T385 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T386 = T387 || mem_valid_received_0;
  assign T387 = memPort_rep_valid && T388;
  assign T388 = memPort_rep_tag == T389;
  assign T389 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T390 = subStateTh_0 == 1'h1/* 1*/;
  assign T391 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T392 = T393 || T257;
  assign T393 = T395 || T394;
  assign T394 = T174 && T5;
  assign T395 = T397 || T396;
  assign T396 = T180 && T5;
  assign T397 = T399 || T398;
  assign T398 = T186 && T5;
  assign T399 = T401 || T400;
  assign T400 = T192 && T5;
  assign T401 = T403 || T402;
  assign T402 = T198 && T5;
  assign T403 = T405 || T404;
  assign T404 = T204 && T5;
  assign T405 = T407 || T406;
  assign T406 = T210 && T5;
  assign T407 = T409 || T408;
  assign T408 = T234 && T5;
  assign T409 = T214 || T410;
  assign T410 = T237 && T22;
  assign T411 = T431 ? 8'hff/* 255*/ : T412;
  assign T412 = T394 ? T430 : T413;
  assign T413 = T396 ? T429 : T414;
  assign T414 = T398 ? T428 : T415;
  assign T415 = T400 ? T427 : T416;
  assign T416 = T402 ? T426 : T417;
  assign T417 = T404 ? T425 : T418;
  assign T418 = T406 ? T424 : T419;
  assign T419 = T408 ? T423 : T420;
  assign T420 = T410 ? T253 : T421;
  assign T421 = T214 ? T422 : State_1;
  assign T422 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T423 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T424 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T425 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T426 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T427 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T428 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T429 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T430 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T431 = T257 || T4;
  assign T432 = subStateTh_1 == 1'h0/* 0*/;
  assign T433 = T435 && T434;
  assign T434 = State_0 == 8'h0/* 0*/;
  assign T435 = subStateTh_0 == 1'h0/* 0*/;
  assign T436 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T437;
  assign T437 = T438[8'ha5/* 165*/:8'h86/* 134*/];
  assign T438 = T582 ? T577 : T439;
  assign T439 = {T576, T575, T574, T573, T440};
  assign T440 = T441[2'h3/* 3*/:1'h0/* 0*/];
  assign T441 = T569 ? T555 : T442;
  assign T442 = {T554, T553, T552, T551, T443};
  assign T443 = T444[2'h3/* 3*/:1'h0/* 0*/];
  assign T444 = T547 ? T542 : T445;
  assign T445 = {T541, T540, T539, T538, T446};
  assign T446 = T447[2'h3/* 3*/:1'h0/* 0*/];
  assign T447 = T534 ? T449 : T448;
  assign T448 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T449 = {memReq4_addr, memReq4_rw, memReq4_cached, memReq4_data, memReq4_size};
  assign memReq4_size = 4'h8/* 8*/;
  assign memReq4_data = T450;
  assign T450 = {64'h0/* 0*/, T451};
  assign T451 = T516 | T452;
  assign T452 = rank_1 & T453;
  assign T453 = {7'h40/* 64*/{T22}};
  assign T454 = T398 || T396;
  assign T455 = T396 ? T496 : T456;
  assign T456 = T398 ? T458 : T457;
  assign T457 = {64'h0/* 0*/, rank_1};
  assign T458 = T487 | T459;
  assign T459 = memRep_1_data & T460;
  assign T460 = {8'h80/* 128*/{T5}};
  assign T461 = T462 || T394;
  assign T462 = T463 || T398;
  assign T463 = T402 || T400;
  assign T464 = T484 ? T465 : memRep_1_data;
  assign T465 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T481 ? T480 : T466;
  assign T466 = {T467};
  assign T467 = T475 | T468;
  assign T468 = memPortReplyStorage_1_data & T469;
  assign T469 = {8'h80/* 128*/{T5}};
  assign T470 = memPort_rep_valid && T471;
  assign T471 = T472[1'h1/* 1*/];
  assign T472 = T473[1'h1/* 1*/:1'h0/* 0*/];
  assign T473 = 2'h1/* 1*/ << memPort_rep_tag;
  assign T474 = T470 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign T475 = memPortReplyStorage_0_data & T476;
  assign T476 = {8'h80/* 128*/{T156}};
  assign T477 = memPort_rep_valid && T478;
  assign T478 = T472[1'h0/* 0*/];
  assign T479 = T477 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T480 = {memPort_rep_bits_data};
  assign T481 = memPort_rep_valid && T482;
  assign T482 = T483 == memPort_rep_tag;
  assign T483 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T484 = T485 || T394;
  assign T485 = T486 || T398;
  assign T486 = T402 || T400;
  assign T487 = memRep_0_data & T488;
  assign T488 = {8'h80/* 128*/{T156}};
  assign T489 = T490 || T173;
  assign T490 = T491 || T185;
  assign T491 = T197 || T191;
  assign T492 = T493 ? T465 : memRep_0_data;
  assign T493 = T494 || T173;
  assign T494 = T495 || T185;
  assign T495 = T197 || T191;
  assign T496 = {64'h0/* 0*/, addOut_out};
  assign addOut_out = T497;
  assign T497 = addPortReplyValue[6'h3f/* 63*/:1'h0/* 0*/];
  assign addPortReplyValue = T513 ? T512 : T498;
  assign T498 = {T499};
  assign T499 = T507 | T500;
  assign T500 = addPortReplyStorage_1_out & T501;
  assign T501 = {7'h40/* 64*/{T5}};
  assign T502 = addPort_rep_valid && T503;
  assign T503 = T504[1'h1/* 1*/];
  assign T504 = T505[1'h1/* 1*/:1'h0/* 0*/];
  assign T505 = 2'h1/* 1*/ << addPort_rep_tag;
  assign T506 = T502 ? addPort_rep_bits_out : addPortReplyStorage_1_out;
  assign addPort_rep_bits_out = mainOff_add_rep_bits_out;
  assign T507 = addPortReplyStorage_0_out & T508;
  assign T508 = {7'h40/* 64*/{T156}};
  assign T509 = addPort_rep_valid && T510;
  assign T510 = T504[1'h0/* 0*/];
  assign T511 = T509 ? addPort_rep_bits_out : addPortReplyStorage_0_out;
  assign T512 = {addPort_rep_bits_out};
  assign T513 = addPort_rep_valid && T514;
  assign T514 = T515 == addPort_rep_tag;
  assign T515 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T516 = rank_0 & T517;
  assign T517 = {7'h40/* 64*/{T76}};
  assign T518 = T185 || T179;
  assign T519 = T179 ? T522 : T520;
  assign T520 = T185 ? T458 : T521;
  assign T521 = {64'h0/* 0*/, rank_0};
  assign T522 = {64'h0/* 0*/, addOut_out};
  assign memReq4_rw = 1'h1/* 1*/;
  assign memReq4_addr = T523;
  assign T523 = T524[5'h1f/* 31*/:1'h0/* 0*/];
  assign T524 = 56'h1000000/* 16777216*/ + T525;
  assign T525 = {21'h0/* 0*/, T526};
  assign T526 = T527 << 32'h3/* 3*/;
  assign T527 = T531 | T528;
  assign T528 = inputReg_1_pageId & T529;
  assign T529 = {6'h20/* 32*/{T22}};
  assign T530 = T214 ? io_in_bits_pageId : inputReg_1_pageId;
  assign T531 = inputReg_0_pageId & T532;
  assign T532 = {6'h20/* 32*/{T76}};
  assign T533 = T225 ? io_in_bits_pageId : inputReg_0_pageId;
  assign T534 = T537 && T535;
  assign T535 = T19 == T536;
  assign T536 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T537 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T538 = T447[8'h83/* 131*/:3'h4/* 4*/];
  assign T539 = T447[8'h84/* 132*/];
  assign T540 = T447[8'h85/* 133*/];
  assign T541 = T447[8'ha5/* 165*/:8'h86/* 134*/];
  assign T542 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h8/* 8*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T543;
  assign T543 = T544[5'h1f/* 31*/:1'h0/* 0*/];
  assign T544 = 56'h1000000/* 16777216*/ + T545;
  assign T545 = {21'h0/* 0*/, T546};
  assign T546 = T527 << 32'h3/* 3*/;
  assign T547 = T550 && T548;
  assign T548 = T19 == T549;
  assign T549 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T550 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T551 = T444[8'h83/* 131*/:3'h4/* 4*/];
  assign T552 = T444[8'h84/* 132*/];
  assign T553 = T444[8'h85/* 133*/];
  assign T554 = T444[8'ha5/* 165*/:8'h86/* 134*/];
  assign T555 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h4/* 4*/;
  assign memReq2_data = T556;
  assign T556 = T560 ^ T557;
  assign T557 = {96'h0/* 0*/, T558};
  assign T558 = 32'h1/* 1*/ << T559;
  assign T559 = T527 & 32'h1f/* 31*/;
  assign T560 = T563 | T561;
  assign T561 = memRep_1_data & T562;
  assign T562 = {8'h80/* 128*/{T22}};
  assign T563 = memRep_0_data & T564;
  assign T564 = {8'h80/* 128*/{T76}};
  assign memReq2_rw = 1'h1/* 1*/;
  assign memReq2_addr = T565;
  assign T565 = T566[5'h1f/* 31*/:1'h0/* 0*/];
  assign T566 = 59'h8000000/* 134217728*/ + T567;
  assign T567 = {27'h0/* 0*/, T568};
  assign T568 = T527 >> 32'h3/* 3*/;
  assign T569 = T572 && T570;
  assign T570 = T19 == T571;
  assign T571 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T572 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T573 = T441[8'h83/* 131*/:3'h4/* 4*/];
  assign T574 = T441[8'h84/* 132*/];
  assign T575 = T441[8'h85/* 133*/];
  assign T576 = T441[8'ha5/* 165*/:8'h86/* 134*/];
  assign T577 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h4/* 4*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T578;
  assign T578 = T579[5'h1f/* 31*/:1'h0/* 0*/];
  assign T579 = 59'h8000000/* 134217728*/ + T580;
  assign T580 = {27'h0/* 0*/, T581};
  assign T581 = T527 >> 32'h3/* 3*/;
  assign T582 = T585 && T583;
  assign T583 = T19 == T584;
  assign T584 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T585 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T586;
  assign T586 = T438[2'h3/* 3*/:1'h0/* 0*/];
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T587;
  assign T587 = T438[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T588;
  assign T588 = T438[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T589;
  assign T589 = T438[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T590;
  assign T590 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mainOff_lock_req_tag = lockPort_req_tag;
  assign lockPort_req_tag = T591;
  assign T591 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign io_out_tag = T592;
  assign T592 = T596 | T593;
  assign T593 = inputTag_1 & T594;
  assign T594 = {4'ha/* 10*/{T22}};
  assign T595 = T214 ? io_in_tag : inputTag_1;
  assign T596 = inputTag_0 & T597;
  assign T597 = {4'ha/* 10*/{T76}};
  assign T598 = T225 ? io_in_tag : inputTag_0;
  RREncode_44 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T147 ),
       .io_valid_1( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T279 ));
  RREncode_45 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T345 ),
       .io_valid_1( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T391 ));
  RREncode_46 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T433 ),
       .io_valid_1( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T436 ));

  always @(posedge clk) begin
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_1 <= T411;
    end
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T26;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T42;
    add_ready_received <= reset ? 1'h0/* 0*/ : T46;
    lock_valid_received_1 <= reset ? 1'h0/* 0*/ : T67;
    lock_valid_received_0 <= reset ? 1'h0/* 0*/ : T77;
    lockPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T87;
    lock_ready_received <= reset ? 1'h0/* 0*/ : T91;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T121;
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T130;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T140;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T144;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T148;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T154) begin
      State_0 <= T241;
    end
    if(T214) begin
      inputReg_1_done <= T223;
    end
    if(T225) begin
      inputReg_0_done <= T227;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T256) begin
      EmitReturnState_1 <= T258;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T262) begin
      EmitReturnState_0 <= T263;
    end
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T287;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    lockPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T318;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T332;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T349;
    lockPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T364;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T378;
    if(T454) begin
      rank_1 <= T455;
    end
    if(T461) begin
      memRep_1_data <= T464;
    end
    if(T470) begin
      memPortReplyStorage_1_data <= T474;
    end
    if(T477) begin
      memPortReplyStorage_0_data <= T479;
    end
    if(T489) begin
      memRep_0_data <= T492;
    end
    if(T502) begin
      addPortReplyStorage_1_out <= T506;
    end
    if(T509) begin
      addPortReplyStorage_0_out <= T511;
    end
    if(T518) begin
      rank_0 <= T519;
    end
    if(T214) begin
      inputReg_1_pageId <= T530;
    end
    if(T225) begin
      inputReg_0_pageId <= T533;
    end
    if(T214) begin
      inputTag_1 <= T595;
    end
    if(T225) begin
      inputTag_0 <= T598;
    end
  end
endmodule

module gPipe_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_5 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_17(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  pcIn0_valid,
    input  pcIn0_bits_request,
    input [15:0] pcIn0_bits_moduleId,
    input [7:0] pcIn0_bits_portId,
    input [19:0] pcIn0_bits_pcValue,
    input [3:0] pcIn0_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag,
    input  io_off_lock_req_ready,
    output io_off_lock_req_valid,
    output[31:0] io_off_lock_req_bits_id,
    output io_off_lock_req_bits_op,
    output[9:0] io_off_lock_req_tag,
    output io_off_lock_rep_ready,
    input  io_off_lock_rep_valid,
    input  io_off_lock_rep_bits_out,
    input [9:0] io_off_lock_rep_tag);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_mainOff_lock_rep_ready;
  wire mainComp_mainOff_lock_req_valid;
  wire mainComp_mainOff_mem_req_valid;
  wire mainComp_io_out_valid;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_mainOff_lock_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_off_lock_rep_ready = mainComp_mainOff_lock_rep_ready;
  assign io_off_lock_req_valid = mainComp_mainOff_lock_req_valid;
  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_off_lock_req_tag = mainComp_mainOff_lock_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateWriter mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_lock_req_ready( io_off_lock_req_ready ),
       .mainOff_lock_req_valid( mainComp_mainOff_lock_req_valid ),
       .mainOff_lock_req_bits_id(  ),
       .mainOff_lock_req_bits_op(  ),
       .mainOff_lock_req_tag( mainComp_mainOff_lock_req_tag ),
       .mainOff_lock_rep_ready( mainComp_mainOff_lock_rep_ready ),
       .mainOff_lock_rep_valid( io_off_lock_rep_valid ),
       .mainOff_lock_rep_bits_out(  ),
       .mainOff_lock_rep_tag( io_off_lock_rep_tag ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_47(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_48(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_49(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateWriter_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_lock_req_ready,
    output mainOff_lock_req_valid,
    output[31:0] mainOff_lock_req_bits_id,
    output mainOff_lock_req_bits_op,
    output[9:0] mainOff_lock_req_tag,
    output mainOff_lock_rep_ready,
    input  mainOff_lock_rep_valid,
    input  mainOff_lock_rep_bits_out,
    input [9:0] mainOff_lock_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire memPort_req_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[4:0] T10;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T11;
  reg[0:0] subStateTh_1;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T15;
  wire AllOffloadsValid_1;
  wire T16;
  wire T17;
  wire T18;
  reg[0:0] addPortHadValidRequest_1;
  wire T19;
  wire T20;
  wire T21;
  wire addPort_req_valid;
  wire T22;
  wire T23;
  wire T24;
  wire[7:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg[0:0] add_valid_received_1;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[9:0] T35;
  wire[9:0] addPort_rep_tag;
  wire addPort_rep_ready;
  wire[9:0] addPort_req_tag;
  wire[9:0] T36;
  wire addPort_rep_valid;
  wire T37;
  wire T38;
  wire[4:0] T39;
  wire T40;
  wire T41;
  reg[0:0] add_valid_received_0;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[9:0] T46;
  wire T47;
  wire T48;
  wire[4:0] T49;
  wire T50;
  wire T51;
  wire[4:0] T52;
  wire T53;
  wire T54;
  wire[4:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[9:0] T59;
  wire T60;
  wire T61;
  wire T62;
  reg[0:0] lockPortHadValidRequest_1;
  wire T63;
  wire T64;
  wire T65;
  wire lockPort_req_valid;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire[7:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  reg[0:0] lock_valid_received_1;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire[9:0] T84;
  wire[9:0] lockPort_rep_tag;
  wire lockPort_rep_valid;
  wire T85;
  wire T86;
  wire[4:0] T87;
  wire T88;
  reg[0:0] lock_valid_received_0;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire[9:0] T93;
  wire T94;
  wire T95;
  wire[4:0] T96;
  wire T97;
  wire T98;
  wire[4:0] T99;
  wire T100;
  wire T101;
  wire[4:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[9:0] T106;
  wire T107;
  wire T108;
  reg[0:0] memPortHadValidRequest_1;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire[4:0] T116;
  wire T117;
  reg[0:0] mem_valid_received_1;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[9:0] T122;
  wire[9:0] memPort_rep_tag;
  wire memPort_rep_valid;
  wire T123;
  wire T124;
  wire[4:0] T125;
  wire T126;
  wire T127;
  wire[9:0] T128;
  wire T129;
  wire T130;
  wire AllOffloadsValid_0;
  wire T131;
  wire T132;
  wire T133;
  reg[0:0] addPortHadValidRequest_0;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] T138;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[9:0] T145;
  wire T146;
  wire T147;
  wire T148;
  reg[0:0] lockPortHadValidRequest_0;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire[4:0] T153;
  wire T154;
  wire T155;
  wire[4:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire[9:0] T160;
  wire T161;
  wire T162;
  reg[0:0] memPortHadValidRequest_0;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire[4:0] T167;
  wire T168;
  wire T169;
  wire[4:0] T170;
  wire T171;
  reg[0:0] mem_valid_received_0;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[9:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire[9:0] T182;
  wire T183;
  reg[0:0] subStateTh_0;
  wire T184;
  wire T185;
  wire T186;
  wire[1:0] T187;
  wire T188;
  wire T189;
  reg[7:0] State_0;
  wire T190;
  wire T191;
  wire T192;
  wire[1:0] T193;
  wire[4:0] T194;
  wire T195;
  wire T196;
  wire[7:0] T197;
  wire[7:0] T198;
  wire[7:0] T199;
  wire[7:0] T200;
  wire T201;
  reg[7:0] State_1;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire[7:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[7:0] T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[7:0] T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[7:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire[7:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[7:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  reg[0:0] inputReg_1_done;
  wire T252;
  wire T253;
  wire[1:0] T254;
  wire[4:0] T255;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire lockPort_rep_ready;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  reg[0:0] inputReg_0_done;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire[7:0] T287;
  wire[7:0] T288;
  wire[7:0] T289;
  wire[7:0] T290;
  wire[7:0] T291;
  wire[7:0] T292;
  wire[7:0] T293;
  wire[7:0] T294;
  wire[7:0] T295;
  wire[7:0] T296;
  wire[7:0] T297;
  wire[7:0] T298;
  wire[7:0] T299;
  wire[7:0] T300;
  wire[7:0] T301;
  reg[7:0] EmitReturnState_1;
  wire T302;
  wire[7:0] T303;
  wire T304;
  wire[7:0] T305;
  wire[7:0] T306;
  reg[7:0] EmitReturnState_0;
  wire T307;
  wire T308;
  wire[7:0] T309;
  wire T310;
  wire[7:0] T311;
  wire[7:0] T312;
  wire[7:0] T313;
  wire[7:0] T314;
  wire[7:0] T315;
  wire[7:0] T316;
  wire[7:0] T317;
  wire[7:0] T318;
  wire T319;
  wire[7:0] T320;
  wire[7:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire[7:0] T342;
  wire[7:0] T343;
  wire[7:0] T344;
  wire[7:0] T345;
  wire[7:0] T346;
  wire[7:0] T347;
  wire[7:0] T348;
  wire[7:0] T349;
  wire[7:0] T350;
  wire[7:0] T351;
  wire[7:0] T352;
  wire[7:0] T353;
  wire[7:0] T354;
  wire[7:0] T355;
  wire[7:0] T356;
  wire[7:0] T357;
  wire[7:0] T358;
  wire[7:0] T359;
  wire[7:0] T360;
  wire[7:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire[1:0] T367;
  wire AllOffloadsReady;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  reg[0:0] addPortHadReadyRequest;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  reg[0:0] add_ready_received;
  wire T377;
  wire T378;
  wire addPort_req_ready;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  reg[0:0] lockPortHadReadyRequest;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  reg[0:0] lock_ready_received;
  wire T389;
  wire T390;
  wire lockPort_req_ready;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  reg[0:0] memPortHadReadyRequest;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  reg[0:0] mem_ready_received;
  wire T400;
  wire T401;
  wire memPort_req_ready;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire[1:0] T411;
  wire T412;
  wire T413;
  wire[7:0] T414;
  wire[7:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[7:0] T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire[7:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T437;
  wire[165:0] T438;
  wire[165:0] T439;
  wire[3:0] T440;
  wire[165:0] T441;
  wire[165:0] T442;
  wire[3:0] T443;
  wire[165:0] T444;
  wire[165:0] T445;
  wire[3:0] T446;
  wire[165:0] T447;
  wire[165:0] T448;
  wire[165:0] T449;
  wire[3:0] memReq4_size;
  wire[127:0] memReq4_data;
  wire[127:0] T450;
  wire[63:0] T451;
  wire[63:0] T452;
  wire[63:0] T453;
  reg[63:0] rank_1;
  wire T454;
  wire[127:0] T455;
  wire[127:0] T456;
  wire[127:0] T457;
  wire[127:0] T458;
  wire[127:0] T459;
  wire[127:0] T460;
  reg[127:0] memRep_1_data;
  wire T461;
  wire T462;
  wire T463;
  wire[127:0] T464;
  wire[127:0] T465;
  wire[127:0] memPortReplyValue;
  wire[127:0] T466;
  wire[127:0] T467;
  wire[127:0] T468;
  wire[127:0] T469;
  reg[127:0] memPortReplyStorage_1_data;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire[1024:0] T473;
  wire[127:0] T474;
  wire[127:0] memPort_rep_bits_data;
  wire[127:0] T475;
  wire[127:0] T476;
  reg[127:0] memPortReplyStorage_0_data;
  wire T477;
  wire T478;
  wire[127:0] T479;
  wire[127:0] T480;
  wire T481;
  wire T482;
  wire[9:0] T483;
  wire T484;
  wire T485;
  wire T486;
  wire[127:0] T487;
  wire[127:0] T488;
  reg[127:0] memRep_0_data;
  wire T489;
  wire T490;
  wire T491;
  wire[127:0] T492;
  wire T493;
  wire T494;
  wire T495;
  wire[127:0] T496;
  wire[63:0] addOut_out;
  wire[63:0] T497;
  wire[63:0] addPortReplyValue;
  wire[63:0] T498;
  wire[63:0] T499;
  wire[63:0] T500;
  wire[63:0] T501;
  reg[63:0] addPortReplyStorage_1_out;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire[1024:0] T505;
  wire[63:0] T506;
  wire[63:0] addPort_rep_bits_out;
  wire[63:0] T507;
  wire[63:0] T508;
  reg[63:0] addPortReplyStorage_0_out;
  wire T509;
  wire T510;
  wire[63:0] T511;
  wire[63:0] T512;
  wire T513;
  wire T514;
  wire[9:0] T515;
  wire[63:0] T516;
  wire[63:0] T517;
  reg[63:0] rank_0;
  wire T518;
  wire[127:0] T519;
  wire[127:0] T520;
  wire[127:0] T521;
  wire[127:0] T522;
  wire memReq4_cached;
  wire memReq4_rw;
  wire[31:0] memReq4_addr;
  wire[31:0] T523;
  wire[55:0] T524;
  wire[55:0] T525;
  wire[34:0] T526;
  wire[31:0] T527;
  wire[31:0] T528;
  wire[31:0] T529;
  reg[31:0] inputReg_1_pageId;
  wire[31:0] T530;
  wire[31:0] T531;
  wire[31:0] T532;
  reg[31:0] inputReg_0_pageId;
  wire[31:0] T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire T537;
  wire[127:0] T538;
  wire T539;
  wire T540;
  wire[31:0] T541;
  wire[165:0] T542;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T543;
  wire[55:0] T544;
  wire[55:0] T545;
  wire[34:0] T546;
  wire T547;
  wire T548;
  wire[7:0] T549;
  wire T550;
  wire[127:0] T551;
  wire T552;
  wire T553;
  wire[31:0] T554;
  wire[165:0] T555;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire[127:0] T556;
  wire[127:0] T557;
  wire[31:0] T558;
  wire[31:0] T559;
  wire[127:0] T560;
  wire[127:0] T561;
  wire[127:0] T562;
  wire[127:0] T563;
  wire[127:0] T564;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T565;
  wire[58:0] T566;
  wire[58:0] T567;
  wire[31:0] T568;
  wire T569;
  wire T570;
  wire[7:0] T571;
  wire T572;
  wire[127:0] T573;
  wire T574;
  wire T575;
  wire[31:0] T576;
  wire[165:0] T577;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T578;
  wire[58:0] T579;
  wire[58:0] T580;
  wire[31:0] T581;
  wire T582;
  wire T583;
  wire[7:0] T584;
  wire T585;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T586;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T587;
  wire memPort_req_bits_cached;
  wire T588;
  wire memPort_req_bits_rw;
  wire T589;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T590;
  wire[9:0] lockPort_req_tag;
  wire[9:0] T591;
  wire[9:0] T592;
  wire[9:0] T593;
  wire[9:0] T594;
  reg[9:0] inputTag_1;
  wire[9:0] T595;
  wire[9:0] T596;
  wire[9:0] T597;
  reg[9:0] inputTag_0;
  wire[9:0] T598;

  assign mainOff_mem_req_valid = memPort_req_valid;
  assign memPort_req_valid = T0;
  assign T0 = T431 && T1;
  assign T1 = T417 || T2;
  assign T2 = T416 && T3;
  assign T3 = T5 == T4;
  assign T4 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T5 = T414 | T6;
  assign T6 = State_1 & T7;
  assign T7 = {4'h8/* 8*/{T8}};
  assign T8 = T9[1'h1/* 1*/];
  assign T9 = T10[1'h1/* 1*/:1'h0/* 0*/];
  assign T10 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T11 = subStateTh_1 == 1'h0/* 0*/;
  assign T12 = T405 ? 1'h1/* 1*/ : T13;
  assign T13 = T14 ? 1'h0/* 0*/ : subStateTh_1;
  assign T14 = T404 == vThreadEncoder_io_chosen;
  assign T15 = T129 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T16;
  assign T16 = T60 && T17;
  assign T17 = T56 || T18;
  assign T18 = ! addPortHadValidRequest_1;
  assign T19 = T53 && T20;
  assign T20 = addPortHadValidRequest_1 || T21;
  assign T21 = T51 && addPort_req_valid;
  assign addPort_req_valid = T22;
  assign T22 = T27 && T23;
  assign T23 = T26 && T24;
  assign T24 = T5 == T25;
  assign T25 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T26 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T27 = T50 && T28;
  assign T28 = ! T29;
  assign T29 = T40 | T30;
  assign T30 = add_valid_received_1 & T8;
  assign T31 = T37 && T32;
  assign T32 = add_valid_received_1 || T33;
  assign T33 = addPort_rep_valid && T34;
  assign T34 = addPort_rep_tag == T35;
  assign T35 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T36;
  assign T36 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T37 = ! T38;
  assign T38 = T39 == 5'h1/* 1*/;
  assign T39 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T40 = add_valid_received_0 & T41;
  assign T41 = T9[1'h0/* 0*/];
  assign T42 = T47 && T43;
  assign T43 = add_valid_received_0 || T44;
  assign T44 = addPort_rep_valid && T45;
  assign T45 = addPort_rep_tag == T46;
  assign T46 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T47 = ! T48;
  assign T48 = T49 == 5'h0/* 0*/;
  assign T49 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T50 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T51 = 5'h1/* 1*/ == T52;
  assign T52 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T53 = ! T54;
  assign T54 = T55 == 5'h1/* 1*/;
  assign T55 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T56 = T57 || add_valid_received_1;
  assign T57 = addPort_rep_valid && T58;
  assign T58 = addPort_rep_tag == T59;
  assign T59 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T60 = T107 && T61;
  assign T61 = T103 || T62;
  assign T62 = ! lockPortHadValidRequest_1;
  assign T63 = T100 && T64;
  assign T64 = lockPortHadValidRequest_1 || T65;
  assign T65 = T98 && lockPort_req_valid;
  assign lockPort_req_valid = T66;
  assign T66 = T76 && T67;
  assign T67 = T72 || T68;
  assign T68 = T71 && T69;
  assign T69 = T5 == T70;
  assign T70 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T72 = T75 && T73;
  assign T73 = T5 == T74;
  assign T74 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T75 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T76 = T97 && T77;
  assign T77 = ! T78;
  assign T78 = T88 | T79;
  assign T79 = lock_valid_received_1 & T8;
  assign T80 = T85 && T81;
  assign T81 = lock_valid_received_1 || T82;
  assign T82 = lockPort_rep_valid && T83;
  assign T83 = lockPort_rep_tag == T84;
  assign T84 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign lockPort_rep_tag = mainOff_lock_rep_tag;
  assign lockPort_rep_valid = mainOff_lock_rep_valid;
  assign T85 = ! T86;
  assign T86 = T87 == 5'h1/* 1*/;
  assign T87 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T88 = lock_valid_received_0 & T41;
  assign T89 = T94 && T90;
  assign T90 = lock_valid_received_0 || T91;
  assign T91 = lockPort_rep_valid && T92;
  assign T92 = lockPort_rep_tag == T93;
  assign T93 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T94 = ! T95;
  assign T95 = T96 == 5'h0/* 0*/;
  assign T96 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T97 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T98 = 5'h1/* 1*/ == T99;
  assign T99 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T100 = ! T101;
  assign T101 = T102 == 5'h1/* 1*/;
  assign T102 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T103 = T104 || lock_valid_received_1;
  assign T104 = lockPort_rep_valid && T105;
  assign T105 = lockPort_rep_tag == T106;
  assign T106 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T107 = T117 || T108;
  assign T108 = ! memPortHadValidRequest_1;
  assign T109 = T114 && T110;
  assign T110 = memPortHadValidRequest_1 || T111;
  assign T111 = T112 && memPort_req_valid;
  assign T112 = 5'h1/* 1*/ == T113;
  assign T113 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T114 = ! T115;
  assign T115 = T116 == 5'h1/* 1*/;
  assign T116 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T117 = T126 || mem_valid_received_1;
  assign T118 = T123 && T119;
  assign T119 = mem_valid_received_1 || T120;
  assign T120 = memPort_rep_valid && T121;
  assign T121 = memPort_rep_tag == T122;
  assign T122 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T123 = ! T124;
  assign T124 = T125 == 5'h1/* 1*/;
  assign T125 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T126 = memPort_rep_valid && T127;
  assign T127 = memPort_rep_tag == T128;
  assign T128 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T129 = subStateTh_1 == 1'h1/* 1*/;
  assign T130 = T183 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T131;
  assign T131 = T146 && T132;
  assign T132 = T142 || T133;
  assign T133 = ! addPortHadValidRequest_0;
  assign T134 = T139 && T135;
  assign T135 = addPortHadValidRequest_0 || T136;
  assign T136 = T137 && addPort_req_valid;
  assign T137 = 5'h0/* 0*/ == T138;
  assign T138 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T139 = ! T140;
  assign T140 = T141 == 5'h0/* 0*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T143 || add_valid_received_0;
  assign T143 = addPort_rep_valid && T144;
  assign T144 = addPort_rep_tag == T145;
  assign T145 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T146 = T161 && T147;
  assign T147 = T157 || T148;
  assign T148 = ! lockPortHadValidRequest_0;
  assign T149 = T154 && T150;
  assign T150 = lockPortHadValidRequest_0 || T151;
  assign T151 = T152 && lockPort_req_valid;
  assign T152 = 5'h0/* 0*/ == T153;
  assign T153 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T154 = ! T155;
  assign T155 = T156 == 5'h0/* 0*/;
  assign T156 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T157 = T158 || lock_valid_received_0;
  assign T158 = lockPort_rep_valid && T159;
  assign T159 = lockPort_rep_tag == T160;
  assign T160 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T161 = T171 || T162;
  assign T162 = ! memPortHadValidRequest_0;
  assign T163 = T168 && T164;
  assign T164 = memPortHadValidRequest_0 || T165;
  assign T165 = T166 && memPort_req_valid;
  assign T166 = 5'h0/* 0*/ == T167;
  assign T167 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T168 = ! T169;
  assign T169 = T170 == 5'h0/* 0*/;
  assign T170 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T171 = T180 || mem_valid_received_0;
  assign T172 = T177 && T173;
  assign T173 = mem_valid_received_0 || T174;
  assign T174 = memPort_rep_valid && T175;
  assign T175 = memPort_rep_tag == T176;
  assign T176 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = memPort_rep_valid && T181;
  assign T181 = memPort_rep_tag == T182;
  assign T182 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T183 = subStateTh_0 == 1'h1/* 1*/;
  assign T184 = T188 ? 1'h1/* 1*/ : T185;
  assign T185 = T186 ? 1'h0/* 0*/ : subStateTh_0;
  assign T186 = T187 == vThreadEncoder_io_chosen;
  assign T187 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T188 = T363 && T189;
  assign T189 = State_0 != 8'hff/* 255*/;
  assign T190 = T323 || T191;
  assign T191 = T195 && T192;
  assign T192 = T193[1'h0/* 0*/];
  assign T193 = T194[1'h1/* 1*/:1'h0/* 0*/];
  assign T194 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T195 = T322 && T196;
  assign T196 = T198 == T197;
  assign T197 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T198 = T320 | T199;
  assign T199 = State_1 & T200;
  assign T200 = {4'h8/* 8*/{T201}};
  assign T201 = T193[1'h1/* 1*/];
  assign T202 = T204 || T203;
  assign T203 = T195 && T201;
  assign T204 = T210 || T205;
  assign T205 = T206 && T201;
  assign T206 = T209 && T207;
  assign T207 = T198 == T208;
  assign T208 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T209 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T210 = T216 || T211;
  assign T211 = T212 && T201;
  assign T212 = T215 && T213;
  assign T213 = T198 == T214;
  assign T214 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T215 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T216 = T222 || T217;
  assign T217 = T218 && T201;
  assign T218 = T221 && T219;
  assign T219 = T198 == T220;
  assign T220 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T221 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T222 = T228 || T223;
  assign T223 = T224 && T201;
  assign T224 = T227 && T225;
  assign T225 = T198 == T226;
  assign T226 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T227 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T228 = T234 || T229;
  assign T229 = T230 && T201;
  assign T230 = T233 && T231;
  assign T231 = T198 == T232;
  assign T232 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T233 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T234 = T240 || T235;
  assign T235 = T236 && T201;
  assign T236 = T239 && T237;
  assign T237 = T198 == T238;
  assign T238 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T239 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T240 = T246 || T241;
  assign T241 = T242 && T201;
  assign T242 = T245 && T243;
  assign T243 = T198 == T244;
  assign T244 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T245 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T246 = T278 || T247;
  assign T247 = T248 && T201;
  assign T248 = T274 && T249;
  assign T249 = ! T250;
  assign T250 = T270 | T251;
  assign T251 = inputReg_1_done & T201;
  assign T252 = T263 && T253;
  assign T253 = T254[1'h1/* 1*/];
  assign T254 = T255[1'h1/* 1*/:1'h0/* 0*/];
  assign T255 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T256 = T258 && T257;
  assign T257 = State_1 == 8'h0/* 0*/;
  assign T258 = subStateTh_1 == 1'h0/* 0*/;
  assign T259 = T261 && T260;
  assign T260 = State_0 == 8'h0/* 0*/;
  assign T261 = subStateTh_0 == 1'h0/* 0*/;
  assign T262 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T263 = T268 && io_in_valid;
  assign mainOff_lock_rep_ready = lockPort_rep_ready;
  assign lockPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_lock_req_valid = lockPort_req_valid;
  assign io_in_ready = T264;
  assign T264 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_valid = T265;
  assign T265 = T267 && T266;
  assign T266 = T5 == 8'hff/* 255*/;
  assign T267 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T268 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T269 = T252 ? io_in_bits_done : inputReg_1_done;
  assign T270 = inputReg_0_done & T192;
  assign T271 = T263 && T272;
  assign T272 = T254[1'h0/* 0*/];
  assign T273 = T271 ? io_in_bits_done : inputReg_0_done;
  assign T274 = T277 && T275;
  assign T275 = T198 == T276;
  assign T276 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T278 = T281 || T279;
  assign T279 = T280 && T201;
  assign T280 = T274 && T250;
  assign T281 = T252 || T282;
  assign T282 = T283 && T8;
  assign T283 = T284 && io_out_ready;
  assign T284 = T286 && T285;
  assign T285 = T5 == 8'hff/* 255*/;
  assign T286 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T287 = T319 ? 8'hff/* 255*/ : T288;
  assign T288 = T211 ? T318 : T289;
  assign T289 = T217 ? T317 : T290;
  assign T290 = T223 ? T316 : T291;
  assign T291 = T229 ? T315 : T292;
  assign T292 = T235 ? T314 : T293;
  assign T293 = T241 ? T313 : T294;
  assign T294 = T247 ? T312 : T295;
  assign T295 = T279 ? T311 : T296;
  assign T296 = T282 ? T299 : T297;
  assign T297 = T252 ? T298 : State_1;
  assign T298 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T299 = T305 | T300;
  assign T300 = EmitReturnState_1 & T301;
  assign T301 = {4'h8/* 8*/{T8}};
  assign T302 = T205 || T203;
  assign T303 = T304 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T304 = T205 || T203;
  assign T305 = EmitReturnState_0 & T306;
  assign T306 = {4'h8/* 8*/{T41}};
  assign T307 = T308 || T191;
  assign T308 = T206 && T192;
  assign T309 = T310 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T310 = T308 || T191;
  assign T311 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T312 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T313 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T314 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T315 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T316 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T317 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T318 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T319 = T205 || T203;
  assign T320 = State_0 & T321;
  assign T321 = {4'h8/* 8*/{T192}};
  assign T322 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T323 = T324 || T308;
  assign T324 = T326 || T325;
  assign T325 = T212 && T192;
  assign T326 = T328 || T327;
  assign T327 = T218 && T192;
  assign T328 = T330 || T329;
  assign T329 = T224 && T192;
  assign T330 = T332 || T331;
  assign T331 = T230 && T192;
  assign T332 = T334 || T333;
  assign T333 = T236 && T192;
  assign T334 = T336 || T335;
  assign T335 = T242 && T192;
  assign T336 = T338 || T337;
  assign T337 = T248 && T192;
  assign T338 = T340 || T339;
  assign T339 = T280 && T192;
  assign T340 = T271 || T341;
  assign T341 = T283 && T41;
  assign T342 = T362 ? 8'hff/* 255*/ : T343;
  assign T343 = T325 ? T361 : T344;
  assign T344 = T327 ? T360 : T345;
  assign T345 = T329 ? T359 : T346;
  assign T346 = T331 ? T358 : T347;
  assign T347 = T333 ? T357 : T348;
  assign T348 = T335 ? T356 : T349;
  assign T349 = T337 ? T355 : T350;
  assign T350 = T339 ? T354 : T351;
  assign T351 = T341 ? T299 : T352;
  assign T352 = T271 ? T353 : State_0;
  assign T353 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T354 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T355 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T356 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T357 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T358 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T359 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T360 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T361 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T362 = T308 || T191;
  assign T363 = T365 && T364;
  assign T364 = State_0 != 8'h0/* 0*/;
  assign T365 = AllOffloadsReady && T366;
  assign T366 = T367 == rThreadEncoder_io_chosen;
  assign T367 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign AllOffloadsReady = T368;
  assign T368 = T380 && T369;
  assign T369 = T376 || T370;
  assign T370 = T372 && T371;
  assign T371 = ! addPort_req_valid;
  assign T372 = ! addPortHadReadyRequest;
  assign T373 = T375 && T374;
  assign T374 = addPortHadReadyRequest || addPort_req_valid;
  assign T375 = ! AllOffloadsReady;
  assign T376 = addPort_req_ready || add_ready_received;
  assign T377 = T379 && T378;
  assign T378 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign T379 = ! AllOffloadsReady;
  assign T380 = T392 && T381;
  assign T381 = T388 || T382;
  assign T382 = T384 && T383;
  assign T383 = ! lockPort_req_valid;
  assign T384 = ! lockPortHadReadyRequest;
  assign T385 = T387 && T386;
  assign T386 = lockPortHadReadyRequest || lockPort_req_valid;
  assign T387 = ! AllOffloadsReady;
  assign T388 = lockPort_req_ready || lock_ready_received;
  assign T389 = T391 && T390;
  assign T390 = lock_ready_received || lockPort_req_ready;
  assign lockPort_req_ready = mainOff_lock_req_ready;
  assign T391 = ! AllOffloadsReady;
  assign T392 = T399 || T393;
  assign T393 = T395 && T394;
  assign T394 = ! memPort_req_valid;
  assign T395 = ! memPortHadReadyRequest;
  assign T396 = T398 && T397;
  assign T397 = memPortHadReadyRequest || memPort_req_valid;
  assign T398 = ! AllOffloadsReady;
  assign T399 = memPort_req_ready || mem_ready_received;
  assign T400 = T402 && T401;
  assign T401 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign T402 = ! AllOffloadsReady;
  assign T403 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T404 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T405 = T407 && T406;
  assign T406 = State_1 != 8'hff/* 255*/;
  assign T407 = T409 && T408;
  assign T408 = State_1 != 8'h0/* 0*/;
  assign T409 = AllOffloadsReady && T410;
  assign T410 = T411 == rThreadEncoder_io_chosen;
  assign T411 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T412 = subStateTh_0 == 1'h0/* 0*/;
  assign T413 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T414 = State_0 & T415;
  assign T415 = {4'h8/* 8*/{T41}};
  assign T416 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T417 = T422 || T418;
  assign T418 = T421 && T419;
  assign T419 = T5 == T420;
  assign T420 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T421 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T422 = T427 || T423;
  assign T423 = T426 && T424;
  assign T424 = T5 == T425;
  assign T425 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T426 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T427 = T430 && T428;
  assign T428 = T5 == T429;
  assign T429 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T430 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T431 = T436 && T432;
  assign T432 = ! T433;
  assign T433 = T435 | T434;
  assign T434 = mem_valid_received_1 & T8;
  assign T435 = mem_valid_received_0 & T41;
  assign T436 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T437;
  assign T437 = T438[8'ha5/* 165*/:8'h86/* 134*/];
  assign T438 = T582 ? T577 : T439;
  assign T439 = {T576, T575, T574, T573, T440};
  assign T440 = T441[2'h3/* 3*/:1'h0/* 0*/];
  assign T441 = T569 ? T555 : T442;
  assign T442 = {T554, T553, T552, T551, T443};
  assign T443 = T444[2'h3/* 3*/:1'h0/* 0*/];
  assign T444 = T547 ? T542 : T445;
  assign T445 = {T541, T540, T539, T538, T446};
  assign T446 = T447[2'h3/* 3*/:1'h0/* 0*/];
  assign T447 = T534 ? T449 : T448;
  assign T448 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T449 = {memReq4_addr, memReq4_rw, memReq4_cached, memReq4_data, memReq4_size};
  assign memReq4_size = 4'h8/* 8*/;
  assign memReq4_data = T450;
  assign T450 = {64'h0/* 0*/, T451};
  assign T451 = T516 | T452;
  assign T452 = rank_1 & T453;
  assign T453 = {7'h40/* 64*/{T8}};
  assign T454 = T223 || T217;
  assign T455 = T217 ? T496 : T456;
  assign T456 = T223 ? T458 : T457;
  assign T457 = {64'h0/* 0*/, rank_1};
  assign T458 = T487 | T459;
  assign T459 = memRep_1_data & T460;
  assign T460 = {8'h80/* 128*/{T201}};
  assign T461 = T462 || T211;
  assign T462 = T463 || T223;
  assign T463 = T235 || T229;
  assign T464 = T484 ? T465 : memRep_1_data;
  assign T465 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T481 ? T480 : T466;
  assign T466 = {T467};
  assign T467 = T475 | T468;
  assign T468 = memPortReplyStorage_1_data & T469;
  assign T469 = {8'h80/* 128*/{T201}};
  assign T470 = memPort_rep_valid && T471;
  assign T471 = T472[1'h1/* 1*/];
  assign T472 = T473[1'h1/* 1*/:1'h0/* 0*/];
  assign T473 = 2'h1/* 1*/ << memPort_rep_tag;
  assign T474 = T470 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign T475 = memPortReplyStorage_0_data & T476;
  assign T476 = {8'h80/* 128*/{T192}};
  assign T477 = memPort_rep_valid && T478;
  assign T478 = T472[1'h0/* 0*/];
  assign T479 = T477 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T480 = {memPort_rep_bits_data};
  assign T481 = memPort_rep_valid && T482;
  assign T482 = T483 == memPort_rep_tag;
  assign T483 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T484 = T485 || T211;
  assign T485 = T486 || T223;
  assign T486 = T235 || T229;
  assign T487 = memRep_0_data & T488;
  assign T488 = {8'h80/* 128*/{T192}};
  assign T489 = T490 || T325;
  assign T490 = T491 || T329;
  assign T491 = T333 || T331;
  assign T492 = T493 ? T465 : memRep_0_data;
  assign T493 = T494 || T325;
  assign T494 = T495 || T329;
  assign T495 = T333 || T331;
  assign T496 = {64'h0/* 0*/, addOut_out};
  assign addOut_out = T497;
  assign T497 = addPortReplyValue[6'h3f/* 63*/:1'h0/* 0*/];
  assign addPortReplyValue = T513 ? T512 : T498;
  assign T498 = {T499};
  assign T499 = T507 | T500;
  assign T500 = addPortReplyStorage_1_out & T501;
  assign T501 = {7'h40/* 64*/{T201}};
  assign T502 = addPort_rep_valid && T503;
  assign T503 = T504[1'h1/* 1*/];
  assign T504 = T505[1'h1/* 1*/:1'h0/* 0*/];
  assign T505 = 2'h1/* 1*/ << addPort_rep_tag;
  assign T506 = T502 ? addPort_rep_bits_out : addPortReplyStorage_1_out;
  assign addPort_rep_bits_out = mainOff_add_rep_bits_out;
  assign T507 = addPortReplyStorage_0_out & T508;
  assign T508 = {7'h40/* 64*/{T192}};
  assign T509 = addPort_rep_valid && T510;
  assign T510 = T504[1'h0/* 0*/];
  assign T511 = T509 ? addPort_rep_bits_out : addPortReplyStorage_0_out;
  assign T512 = {addPort_rep_bits_out};
  assign T513 = addPort_rep_valid && T514;
  assign T514 = T515 == addPort_rep_tag;
  assign T515 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T516 = rank_0 & T517;
  assign T517 = {7'h40/* 64*/{T41}};
  assign T518 = T329 || T327;
  assign T519 = T327 ? T522 : T520;
  assign T520 = T329 ? T458 : T521;
  assign T521 = {64'h0/* 0*/, rank_0};
  assign T522 = {64'h0/* 0*/, addOut_out};
  assign memReq4_rw = 1'h1/* 1*/;
  assign memReq4_addr = T523;
  assign T523 = T524[5'h1f/* 31*/:1'h0/* 0*/];
  assign T524 = 56'h1000000/* 16777216*/ + T525;
  assign T525 = {21'h0/* 0*/, T526};
  assign T526 = T527 << 32'h3/* 3*/;
  assign T527 = T531 | T528;
  assign T528 = inputReg_1_pageId & T529;
  assign T529 = {6'h20/* 32*/{T8}};
  assign T530 = T252 ? io_in_bits_pageId : inputReg_1_pageId;
  assign T531 = inputReg_0_pageId & T532;
  assign T532 = {6'h20/* 32*/{T41}};
  assign T533 = T271 ? io_in_bits_pageId : inputReg_0_pageId;
  assign T534 = T537 && T535;
  assign T535 = T5 == T536;
  assign T536 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T537 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T538 = T447[8'h83/* 131*/:3'h4/* 4*/];
  assign T539 = T447[8'h84/* 132*/];
  assign T540 = T447[8'h85/* 133*/];
  assign T541 = T447[8'ha5/* 165*/:8'h86/* 134*/];
  assign T542 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h8/* 8*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T543;
  assign T543 = T544[5'h1f/* 31*/:1'h0/* 0*/];
  assign T544 = 56'h1000000/* 16777216*/ + T545;
  assign T545 = {21'h0/* 0*/, T546};
  assign T546 = T527 << 32'h3/* 3*/;
  assign T547 = T550 && T548;
  assign T548 = T5 == T549;
  assign T549 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T550 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T551 = T444[8'h83/* 131*/:3'h4/* 4*/];
  assign T552 = T444[8'h84/* 132*/];
  assign T553 = T444[8'h85/* 133*/];
  assign T554 = T444[8'ha5/* 165*/:8'h86/* 134*/];
  assign T555 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h4/* 4*/;
  assign memReq2_data = T556;
  assign T556 = T560 ^ T557;
  assign T557 = {96'h0/* 0*/, T558};
  assign T558 = 32'h1/* 1*/ << T559;
  assign T559 = T527 & 32'h1f/* 31*/;
  assign T560 = T563 | T561;
  assign T561 = memRep_1_data & T562;
  assign T562 = {8'h80/* 128*/{T8}};
  assign T563 = memRep_0_data & T564;
  assign T564 = {8'h80/* 128*/{T41}};
  assign memReq2_rw = 1'h1/* 1*/;
  assign memReq2_addr = T565;
  assign T565 = T566[5'h1f/* 31*/:1'h0/* 0*/];
  assign T566 = 59'h8000000/* 134217728*/ + T567;
  assign T567 = {27'h0/* 0*/, T568};
  assign T568 = T527 >> 32'h3/* 3*/;
  assign T569 = T572 && T570;
  assign T570 = T5 == T571;
  assign T571 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T572 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T573 = T441[8'h83/* 131*/:3'h4/* 4*/];
  assign T574 = T441[8'h84/* 132*/];
  assign T575 = T441[8'h85/* 133*/];
  assign T576 = T441[8'ha5/* 165*/:8'h86/* 134*/];
  assign T577 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h4/* 4*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T578;
  assign T578 = T579[5'h1f/* 31*/:1'h0/* 0*/];
  assign T579 = 59'h8000000/* 134217728*/ + T580;
  assign T580 = {27'h0/* 0*/, T581};
  assign T581 = T527 >> 32'h3/* 3*/;
  assign T582 = T585 && T583;
  assign T583 = T5 == T584;
  assign T584 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T585 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T586;
  assign T586 = T438[2'h3/* 3*/:1'h0/* 0*/];
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T587;
  assign T587 = T438[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T588;
  assign T588 = T438[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T589;
  assign T589 = T438[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T590;
  assign T590 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mainOff_lock_req_tag = lockPort_req_tag;
  assign lockPort_req_tag = T591;
  assign T591 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign io_out_tag = T592;
  assign T592 = T596 | T593;
  assign T593 = inputTag_1 & T594;
  assign T594 = {4'ha/* 10*/{T8}};
  assign T595 = T252 ? io_in_tag : inputTag_1;
  assign T596 = inputTag_0 & T597;
  assign T597 = {4'ha/* 10*/{T41}};
  assign T598 = T271 ? io_in_tag : inputTag_0;
  RREncode_47 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T412 ),
       .io_valid_1( T11 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T413 ));
  RREncode_48 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T130 ),
       .io_valid_1( T15 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T403 ));
  RREncode_49 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T259 ),
       .io_valid_1( T256 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T262 ));

  always @(posedge clk) begin
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T12;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T19;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T31;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T42;
    lockPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T63;
    lock_valid_received_1 <= reset ? 1'h0/* 0*/ : T80;
    lock_valid_received_0 <= reset ? 1'h0/* 0*/ : T89;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T109;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T118;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T134;
    lockPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T149;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T163;
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T172;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T184;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T190) begin
      State_0 <= T342;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T202) begin
      State_1 <= T287;
    end
    if(T252) begin
      inputReg_1_done <= T269;
    end
    if(T271) begin
      inputReg_0_done <= T273;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T302) begin
      EmitReturnState_1 <= T303;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T307) begin
      EmitReturnState_0 <= T309;
    end
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T373;
    add_ready_received <= reset ? 1'h0/* 0*/ : T377;
    lockPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T385;
    lock_ready_received <= reset ? 1'h0/* 0*/ : T389;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T396;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T400;
    if(T454) begin
      rank_1 <= T455;
    end
    if(T461) begin
      memRep_1_data <= T464;
    end
    if(T470) begin
      memPortReplyStorage_1_data <= T474;
    end
    if(T477) begin
      memPortReplyStorage_0_data <= T479;
    end
    if(T489) begin
      memRep_0_data <= T492;
    end
    if(T502) begin
      addPortReplyStorage_1_out <= T506;
    end
    if(T509) begin
      addPortReplyStorage_0_out <= T511;
    end
    if(T518) begin
      rank_0 <= T519;
    end
    if(T252) begin
      inputReg_1_pageId <= T530;
    end
    if(T271) begin
      inputReg_0_pageId <= T533;
    end
    if(T252) begin
      inputTag_1 <= T595;
    end
    if(T271) begin
      inputTag_0 <= T598;
    end
  end
endmodule

module gPipe_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_6 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_18(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag,
    input  io_off_lock_req_ready,
    output io_off_lock_req_valid,
    output[31:0] io_off_lock_req_bits_id,
    output io_off_lock_req_bits_op,
    output[9:0] io_off_lock_req_tag,
    output io_off_lock_rep_ready,
    input  io_off_lock_rep_valid,
    input  io_off_lock_rep_bits_out,
    input [9:0] io_off_lock_rep_tag);

  wire mainComp_mainOff_mem_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire mainComp_mainOff_lock_rep_ready;
  wire mainComp_mainOff_lock_req_valid;
  wire mainComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_mainOff_lock_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_off_lock_rep_ready = mainComp_mainOff_lock_rep_ready;
  assign io_off_lock_req_valid = mainComp_mainOff_lock_req_valid;
  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_off_lock_req_tag = mainComp_mainOff_lock_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateWriter_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_lock_req_ready( io_off_lock_req_ready ),
       .mainOff_lock_req_valid( mainComp_mainOff_lock_req_valid ),
       .mainOff_lock_req_bits_id(  ),
       .mainOff_lock_req_bits_op(  ),
       .mainOff_lock_req_tag( mainComp_mainOff_lock_req_tag ),
       .mainOff_lock_rep_ready( mainComp_mainOff_lock_rep_ready ),
       .mainOff_lock_rep_valid( io_off_lock_rep_valid ),
       .mainOff_lock_rep_bits_out(  ),
       .mainOff_lock_rep_tag( io_off_lock_rep_tag ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_5 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_50(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_51(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_52(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateWriter_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_lock_req_ready,
    output mainOff_lock_req_valid,
    output[31:0] mainOff_lock_req_bits_id,
    output mainOff_lock_req_bits_op,
    output[9:0] mainOff_lock_req_tag,
    output mainOff_lock_rep_ready,
    input  mainOff_lock_rep_valid,
    input  mainOff_lock_rep_bits_out,
    input [9:0] mainOff_lock_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire lockPort_req_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[7:0] T4;
  wire[7:0] T5;
  wire[7:0] T6;
  wire[7:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[4:0] T10;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T11;
  reg[0:0] subStateTh_1;
  wire T12;
  wire T13;
  wire T14;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T15;
  wire AllOffloadsValid_1;
  wire T16;
  wire T17;
  wire T18;
  reg[0:0] addPortHadValidRequest_1;
  wire T19;
  wire T20;
  wire T21;
  wire addPort_req_valid;
  wire T22;
  wire T23;
  wire T24;
  wire[7:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg[0:0] add_valid_received_1;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[9:0] T35;
  wire[9:0] addPort_rep_tag;
  wire addPort_rep_ready;
  wire[9:0] addPort_req_tag;
  wire[9:0] T36;
  wire addPort_rep_valid;
  wire T37;
  wire T38;
  wire[4:0] T39;
  wire T40;
  wire T41;
  reg[0:0] add_valid_received_0;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[9:0] T46;
  wire T47;
  wire T48;
  wire[4:0] T49;
  wire T50;
  wire T51;
  wire[4:0] T52;
  wire T53;
  wire T54;
  wire[4:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire[9:0] T59;
  wire T60;
  wire T61;
  wire T62;
  reg[0:0] lockPortHadValidRequest_1;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[4:0] T67;
  wire T68;
  wire T69;
  wire[4:0] T70;
  wire T71;
  reg[0:0] lock_valid_received_1;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[9:0] T76;
  wire[9:0] lockPort_rep_tag;
  wire lockPort_rep_valid;
  wire T77;
  wire T78;
  wire[4:0] T79;
  wire T80;
  wire T81;
  wire[9:0] T82;
  wire T83;
  wire T84;
  reg[0:0] memPortHadValidRequest_1;
  wire T85;
  wire T86;
  wire T87;
  wire memPort_req_valid;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[7:0] T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[7:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[7:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] mem_valid_received_1;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[9:0] T116;
  wire[9:0] memPort_rep_tag;
  wire lockPort_rep_ready;
  wire T117;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T118;
  wire T119;
  reg[7:0] State_1;
  wire T120;
  wire T121;
  wire T122;
  wire[1:0] T123;
  wire[4:0] T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire[7:0] T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[7:0] T131;
  wire[7:0] T132;
  wire T133;
  reg[7:0] State_0;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[7:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire[7:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[7:0] T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire[7:0] T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[7:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[7:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  reg[0:0] inputReg_1_done;
  wire T184;
  wire T185;
  wire[1:0] T186;
  wire[4:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg[0:0] inputReg_0_done;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[7:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire[7:0] T211;
  wire[7:0] T212;
  wire[7:0] T213;
  wire[7:0] T214;
  wire[7:0] T215;
  wire[7:0] T216;
  wire[7:0] T217;
  wire[7:0] T218;
  wire[7:0] T219;
  wire[7:0] T220;
  wire[7:0] T221;
  wire[7:0] T222;
  wire[7:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  reg[7:0] EmitReturnState_1;
  wire T226;
  wire T227;
  wire[7:0] T228;
  wire T229;
  wire[7:0] T230;
  wire[7:0] T231;
  reg[7:0] EmitReturnState_0;
  wire T232;
  wire[7:0] T233;
  wire T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire[7:0] T240;
  wire[7:0] T241;
  wire[7:0] T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[7:0] T266;
  wire[7:0] T267;
  wire[7:0] T268;
  wire[7:0] T269;
  wire[7:0] T270;
  wire[7:0] T271;
  wire[7:0] T272;
  wire[7:0] T273;
  wire[7:0] T274;
  wire[7:0] T275;
  wire[7:0] T276;
  wire[7:0] T277;
  wire[7:0] T278;
  wire[7:0] T279;
  wire[7:0] T280;
  wire[7:0] T281;
  wire[7:0] T282;
  wire[7:0] T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  reg[0:0] subStateTh_0;
  wire T289;
  wire T290;
  wire T291;
  wire[1:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire[1:0] T299;
  wire AllOffloadsReady;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  reg[0:0] addPortHadReadyRequest;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  reg[0:0] add_ready_received;
  wire T309;
  wire T310;
  wire addPort_req_ready;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  reg[0:0] lockPortHadReadyRequest;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  reg[0:0] lock_ready_received;
  wire T321;
  wire T322;
  wire lockPort_req_ready;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  reg[0:0] memPortHadReadyRequest;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  reg[0:0] mem_ready_received;
  wire T332;
  wire T333;
  wire memPort_req_ready;
  wire T334;
  wire T335;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T336;
  wire[165:0] T337;
  wire[165:0] T338;
  wire[3:0] T339;
  wire[165:0] T340;
  wire[165:0] T341;
  wire[3:0] T342;
  wire[165:0] T343;
  wire[165:0] T344;
  wire[3:0] T345;
  wire[165:0] T346;
  wire[165:0] T347;
  wire[165:0] T348;
  wire[3:0] memReq4_size;
  wire[127:0] memReq4_data;
  wire[127:0] T349;
  wire[63:0] T350;
  wire[63:0] T351;
  wire[63:0] T352;
  reg[63:0] rank_1;
  wire T353;
  wire[127:0] T354;
  wire[127:0] T355;
  wire[127:0] T356;
  wire[127:0] T357;
  wire[127:0] T358;
  wire[127:0] T359;
  reg[127:0] memRep_1_data;
  wire T360;
  wire T361;
  wire T362;
  wire[127:0] T363;
  wire[127:0] T364;
  wire[127:0] memPortReplyValue;
  wire[127:0] T365;
  wire[127:0] T366;
  wire[127:0] T367;
  wire[127:0] T368;
  reg[127:0] memPortReplyStorage_1_data;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1024:0] T372;
  wire memPort_rep_valid;
  wire[127:0] T373;
  wire[127:0] memPort_rep_bits_data;
  wire[127:0] T374;
  wire[127:0] T375;
  reg[127:0] memPortReplyStorage_0_data;
  wire T376;
  wire T377;
  wire[127:0] T378;
  wire[127:0] T379;
  wire T380;
  wire T381;
  wire[9:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire[127:0] T386;
  wire[127:0] T387;
  reg[127:0] memRep_0_data;
  wire T388;
  wire T389;
  wire T390;
  wire[127:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[127:0] T395;
  wire[63:0] addOut_out;
  wire[63:0] T396;
  wire[63:0] addPortReplyValue;
  wire[63:0] T397;
  wire[63:0] T398;
  wire[63:0] T399;
  wire[63:0] T400;
  reg[63:0] addPortReplyStorage_1_out;
  wire T401;
  wire T402;
  wire[1:0] T403;
  wire[1024:0] T404;
  wire[63:0] T405;
  wire[63:0] addPort_rep_bits_out;
  wire[63:0] T406;
  wire[63:0] T407;
  reg[63:0] addPortReplyStorage_0_out;
  wire T408;
  wire T409;
  wire[63:0] T410;
  wire[63:0] T411;
  wire T412;
  wire T413;
  wire[9:0] T414;
  wire[63:0] T415;
  wire[63:0] T416;
  reg[63:0] rank_0;
  wire T417;
  wire[127:0] T418;
  wire[127:0] T419;
  wire[127:0] T420;
  wire[127:0] T421;
  wire memReq4_cached;
  wire memReq4_rw;
  wire[31:0] memReq4_addr;
  wire[31:0] T422;
  wire[55:0] T423;
  wire[55:0] T424;
  wire[34:0] T425;
  wire[31:0] T426;
  wire[31:0] T427;
  wire[31:0] T428;
  reg[31:0] inputReg_1_pageId;
  wire[31:0] T429;
  wire[31:0] T430;
  wire[31:0] T431;
  reg[31:0] inputReg_0_pageId;
  wire[31:0] T432;
  wire T433;
  wire T434;
  wire[7:0] T435;
  wire T436;
  wire[127:0] T437;
  wire T438;
  wire T439;
  wire[31:0] T440;
  wire[165:0] T441;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T442;
  wire[55:0] T443;
  wire[55:0] T444;
  wire[34:0] T445;
  wire T446;
  wire T447;
  wire[7:0] T448;
  wire T449;
  wire[127:0] T450;
  wire T451;
  wire T452;
  wire[31:0] T453;
  wire[165:0] T454;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire[127:0] T455;
  wire[127:0] T456;
  wire[31:0] T457;
  wire[31:0] T458;
  wire[127:0] T459;
  wire[127:0] T460;
  wire[127:0] T461;
  wire[127:0] T462;
  wire[127:0] T463;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T464;
  wire[58:0] T465;
  wire[58:0] T466;
  wire[31:0] T467;
  wire T468;
  wire T469;
  wire[7:0] T470;
  wire T471;
  wire[127:0] T472;
  wire T473;
  wire T474;
  wire[31:0] T475;
  wire[165:0] T476;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T477;
  wire[58:0] T478;
  wire[58:0] T479;
  wire[31:0] T480;
  wire T481;
  wire T482;
  wire[7:0] T483;
  wire T484;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T485;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T486;
  wire memPort_req_bits_cached;
  wire T487;
  wire memPort_req_bits_rw;
  wire T488;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T489;
  wire T490;
  wire T491;
  wire[4:0] T492;
  wire T493;
  reg[0:0] mem_valid_received_0;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire[9:0] T498;
  wire T499;
  wire T500;
  wire[4:0] T501;
  wire T502;
  wire T503;
  wire[4:0] T504;
  wire T505;
  wire T506;
  wire[4:0] T507;
  wire T508;
  wire T509;
  wire T510;
  wire[9:0] T511;
  wire T512;
  wire T513;
  wire AllOffloadsValid_0;
  wire T514;
  wire T515;
  wire T516;
  reg[0:0] addPortHadValidRequest_0;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire[4:0] T521;
  wire T522;
  wire T523;
  wire[4:0] T524;
  wire T525;
  wire T526;
  wire T527;
  wire[9:0] T528;
  wire T529;
  wire T530;
  wire T531;
  reg[0:0] lockPortHadValidRequest_0;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[4:0] T536;
  wire T537;
  wire T538;
  wire[4:0] T539;
  wire T540;
  reg[0:0] lock_valid_received_0;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire[9:0] T545;
  wire T546;
  wire T547;
  wire[4:0] T548;
  wire T549;
  wire T550;
  wire[9:0] T551;
  wire T552;
  wire T553;
  reg[0:0] memPortHadValidRequest_0;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[4:0] T558;
  wire T559;
  wire T560;
  wire[4:0] T561;
  wire T562;
  wire T563;
  wire T564;
  wire[9:0] T565;
  wire T566;
  wire T567;
  wire[1:0] T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire[1:0] T575;
  wire T576;
  wire T577;
  wire[7:0] T578;
  wire[7:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire[7:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire[9:0] lockPort_req_tag;
  wire[9:0] T591;
  wire[9:0] T592;
  wire[9:0] T593;
  wire[9:0] T594;
  reg[9:0] inputTag_1;
  wire[9:0] T595;
  wire[9:0] T596;
  wire[9:0] T597;
  reg[9:0] inputTag_0;
  wire[9:0] T598;

  assign mainOff_lock_req_valid = lockPort_req_valid;
  assign lockPort_req_valid = T0;
  assign T0 = T585 && T1;
  assign T1 = T581 || T2;
  assign T2 = T580 && T3;
  assign T3 = T5 == T4;
  assign T4 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T5 = T578 | T6;
  assign T6 = State_1 & T7;
  assign T7 = {4'h8/* 8*/{T8}};
  assign T8 = T9[1'h1/* 1*/];
  assign T9 = T10[1'h1/* 1*/:1'h0/* 0*/];
  assign T10 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T11 = subStateTh_1 == 1'h0/* 0*/;
  assign T12 = T569 ? 1'h1/* 1*/ : T13;
  assign T13 = T14 ? 1'h0/* 0*/ : subStateTh_1;
  assign T14 = T568 == vThreadEncoder_io_chosen;
  assign T15 = T512 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T16;
  assign T16 = T60 && T17;
  assign T17 = T56 || T18;
  assign T18 = ! addPortHadValidRequest_1;
  assign T19 = T53 && T20;
  assign T20 = addPortHadValidRequest_1 || T21;
  assign T21 = T51 && addPort_req_valid;
  assign addPort_req_valid = T22;
  assign T22 = T27 && T23;
  assign T23 = T26 && T24;
  assign T24 = T5 == T25;
  assign T25 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T26 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T27 = T50 && T28;
  assign T28 = ! T29;
  assign T29 = T40 | T30;
  assign T30 = add_valid_received_1 & T8;
  assign T31 = T37 && T32;
  assign T32 = add_valid_received_1 || T33;
  assign T33 = addPort_rep_valid && T34;
  assign T34 = addPort_rep_tag == T35;
  assign T35 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T36;
  assign T36 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T37 = ! T38;
  assign T38 = T39 == 5'h1/* 1*/;
  assign T39 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T40 = add_valid_received_0 & T41;
  assign T41 = T9[1'h0/* 0*/];
  assign T42 = T47 && T43;
  assign T43 = add_valid_received_0 || T44;
  assign T44 = addPort_rep_valid && T45;
  assign T45 = addPort_rep_tag == T46;
  assign T46 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T47 = ! T48;
  assign T48 = T49 == 5'h0/* 0*/;
  assign T49 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T50 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T51 = 5'h1/* 1*/ == T52;
  assign T52 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T53 = ! T54;
  assign T54 = T55 == 5'h1/* 1*/;
  assign T55 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T56 = T57 || add_valid_received_1;
  assign T57 = addPort_rep_valid && T58;
  assign T58 = addPort_rep_tag == T59;
  assign T59 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T60 = T83 && T61;
  assign T61 = T71 || T62;
  assign T62 = ! lockPortHadValidRequest_1;
  assign T63 = T68 && T64;
  assign T64 = lockPortHadValidRequest_1 || T65;
  assign T65 = T66 && lockPort_req_valid;
  assign T66 = 5'h1/* 1*/ == T67;
  assign T67 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T68 = ! T69;
  assign T69 = T70 == 5'h1/* 1*/;
  assign T70 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T71 = T80 || lock_valid_received_1;
  assign T72 = T77 && T73;
  assign T73 = lock_valid_received_1 || T74;
  assign T74 = lockPort_rep_valid && T75;
  assign T75 = lockPort_rep_tag == T76;
  assign T76 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign lockPort_rep_tag = mainOff_lock_rep_tag;
  assign lockPort_rep_valid = mainOff_lock_rep_valid;
  assign T77 = ! T78;
  assign T78 = T79 == 5'h1/* 1*/;
  assign T79 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T80 = lockPort_rep_valid && T81;
  assign T81 = lockPort_rep_tag == T82;
  assign T82 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T83 = T508 || T84;
  assign T84 = ! memPortHadValidRequest_1;
  assign T85 = T505 && T86;
  assign T86 = memPortHadValidRequest_1 || T87;
  assign T87 = T503 && memPort_req_valid;
  assign memPort_req_valid = T88;
  assign T88 = T108 && T89;
  assign T89 = T94 || T90;
  assign T90 = T93 && T91;
  assign T91 = T5 == T92;
  assign T92 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T93 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T94 = T99 || T95;
  assign T95 = T98 && T96;
  assign T96 = T5 == T97;
  assign T97 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T98 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T99 = T104 || T100;
  assign T100 = T103 && T101;
  assign T101 = T5 == T102;
  assign T102 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T103 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T104 = T107 && T105;
  assign T105 = T5 == T106;
  assign T106 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T107 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T108 = T502 && T109;
  assign T109 = ! T110;
  assign T110 = T493 | T111;
  assign T111 = mem_valid_received_1 & T8;
  assign T112 = T490 && T113;
  assign T113 = mem_valid_received_1 || T114;
  assign T114 = memPort_rep_valid && T115;
  assign T115 = memPort_rep_tag == T116;
  assign T116 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign mainOff_mem_req_valid = memPort_req_valid;
  assign mainOff_lock_rep_ready = lockPort_rep_ready;
  assign lockPort_rep_ready = 1'h1/* 1*/;
  assign io_in_ready = T117;
  assign T117 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T118 = T285 && T119;
  assign T119 = State_1 == 8'h0/* 0*/;
  assign T120 = T245 || T121;
  assign T121 = T125 && T122;
  assign T122 = T123[1'h1/* 1*/];
  assign T123 = T124[1'h1/* 1*/:1'h0/* 0*/];
  assign T124 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T125 = T244 && T126;
  assign T126 = T128 == T127;
  assign T127 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T128 = T131 | T129;
  assign T129 = State_1 & T130;
  assign T130 = {4'h8/* 8*/{T122}};
  assign T131 = State_0 & T132;
  assign T132 = {4'h8/* 8*/{T133}};
  assign T133 = T123[1'h0/* 0*/];
  assign T134 = T136 || T135;
  assign T135 = T125 && T133;
  assign T136 = T142 || T137;
  assign T137 = T138 && T133;
  assign T138 = T141 && T139;
  assign T139 = T128 == T140;
  assign T140 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T141 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T142 = T148 || T143;
  assign T143 = T144 && T133;
  assign T144 = T147 && T145;
  assign T145 = T128 == T146;
  assign T146 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T147 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T148 = T154 || T149;
  assign T149 = T150 && T133;
  assign T150 = T153 && T151;
  assign T151 = T128 == T152;
  assign T152 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T153 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T154 = T160 || T155;
  assign T155 = T156 && T133;
  assign T156 = T159 && T157;
  assign T157 = T128 == T158;
  assign T158 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T159 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T160 = T166 || T161;
  assign T161 = T162 && T133;
  assign T162 = T165 && T163;
  assign T163 = T128 == T164;
  assign T164 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T165 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T166 = T172 || T167;
  assign T167 = T168 && T133;
  assign T168 = T171 && T169;
  assign T169 = T128 == T170;
  assign T170 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T171 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T172 = T178 || T173;
  assign T173 = T174 && T133;
  assign T174 = T177 && T175;
  assign T175 = T128 == T176;
  assign T176 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T177 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T178 = T199 || T179;
  assign T179 = T180 && T133;
  assign T180 = T195 && T181;
  assign T181 = ! T182;
  assign T182 = T191 | T183;
  assign T183 = inputReg_1_done & T122;
  assign T184 = T188 && T185;
  assign T185 = T186[1'h1/* 1*/];
  assign T186 = T187[1'h1/* 1*/:1'h0/* 0*/];
  assign T187 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T188 = T189 && io_in_valid;
  assign T189 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T190 = T184 ? io_in_bits_done : inputReg_1_done;
  assign T191 = inputReg_0_done & T133;
  assign T192 = T188 && T193;
  assign T193 = T186[1'h0/* 0*/];
  assign T194 = T192 ? io_in_bits_done : inputReg_0_done;
  assign T195 = T198 && T196;
  assign T196 = T128 == T197;
  assign T197 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T198 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T199 = T202 || T200;
  assign T200 = T201 && T133;
  assign T201 = T195 && T182;
  assign T202 = T192 || T203;
  assign T203 = T204 && T41;
  assign T204 = T208 && io_out_ready;
  assign io_out_valid = T205;
  assign T205 = T207 && T206;
  assign T206 = T5 == 8'hff/* 255*/;
  assign T207 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T208 = T210 && T209;
  assign T209 = T5 == 8'hff/* 255*/;
  assign T210 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T211 = T243 ? 8'hff/* 255*/ : T212;
  assign T212 = T143 ? T242 : T213;
  assign T213 = T149 ? T241 : T214;
  assign T214 = T155 ? T240 : T215;
  assign T215 = T161 ? T239 : T216;
  assign T216 = T167 ? T238 : T217;
  assign T217 = T173 ? T237 : T218;
  assign T218 = T179 ? T236 : T219;
  assign T219 = T200 ? T235 : T220;
  assign T220 = T203 ? T223 : T221;
  assign T221 = T192 ? T222 : State_0;
  assign T222 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T223 = T230 | T224;
  assign T224 = EmitReturnState_1 & T225;
  assign T225 = {4'h8/* 8*/{T8}};
  assign T226 = T227 || T121;
  assign T227 = T138 && T122;
  assign T228 = T229 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T229 = T227 || T121;
  assign T230 = EmitReturnState_0 & T231;
  assign T231 = {4'h8/* 8*/{T41}};
  assign T232 = T137 || T135;
  assign T233 = T234 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T234 = T137 || T135;
  assign T235 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T236 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T237 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T238 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T239 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T240 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T241 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T242 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T243 = T137 || T135;
  assign T244 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T245 = T246 || T227;
  assign T246 = T248 || T247;
  assign T247 = T144 && T122;
  assign T248 = T250 || T249;
  assign T249 = T150 && T122;
  assign T250 = T252 || T251;
  assign T251 = T156 && T122;
  assign T252 = T254 || T253;
  assign T253 = T162 && T122;
  assign T254 = T256 || T255;
  assign T255 = T168 && T122;
  assign T256 = T258 || T257;
  assign T257 = T174 && T122;
  assign T258 = T260 || T259;
  assign T259 = T180 && T122;
  assign T260 = T262 || T261;
  assign T261 = T201 && T122;
  assign T262 = T184 || T263;
  assign T263 = T204 && T8;
  assign T264 = T284 ? 8'hff/* 255*/ : T265;
  assign T265 = T247 ? T283 : T266;
  assign T266 = T249 ? T282 : T267;
  assign T267 = T251 ? T281 : T268;
  assign T268 = T253 ? T280 : T269;
  assign T269 = T255 ? T279 : T270;
  assign T270 = T257 ? T278 : T271;
  assign T271 = T259 ? T277 : T272;
  assign T272 = T261 ? T276 : T273;
  assign T273 = T263 ? T223 : T274;
  assign T274 = T184 ? T275 : State_1;
  assign T275 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T276 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T277 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T278 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T279 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T280 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T281 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T282 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T283 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T284 = T227 || T121;
  assign T285 = subStateTh_1 == 1'h0/* 0*/;
  assign T286 = T288 && T287;
  assign T287 = State_0 == 8'h0/* 0*/;
  assign T288 = subStateTh_0 == 1'h0/* 0*/;
  assign T289 = T293 ? 1'h1/* 1*/ : T290;
  assign T290 = T291 ? 1'h0/* 0*/ : subStateTh_0;
  assign T291 = T292 == vThreadEncoder_io_chosen;
  assign T292 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T293 = T295 && T294;
  assign T294 = State_0 != 8'hff/* 255*/;
  assign T295 = T297 && T296;
  assign T296 = State_0 != 8'h0/* 0*/;
  assign T297 = AllOffloadsReady && T298;
  assign T298 = T299 == rThreadEncoder_io_chosen;
  assign T299 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign AllOffloadsReady = T300;
  assign T300 = T312 && T301;
  assign T301 = T308 || T302;
  assign T302 = T304 && T303;
  assign T303 = ! addPort_req_valid;
  assign T304 = ! addPortHadReadyRequest;
  assign T305 = T307 && T306;
  assign T306 = addPortHadReadyRequest || addPort_req_valid;
  assign T307 = ! AllOffloadsReady;
  assign T308 = addPort_req_ready || add_ready_received;
  assign T309 = T311 && T310;
  assign T310 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign T311 = ! AllOffloadsReady;
  assign T312 = T324 && T313;
  assign T313 = T320 || T314;
  assign T314 = T316 && T315;
  assign T315 = ! lockPort_req_valid;
  assign T316 = ! lockPortHadReadyRequest;
  assign T317 = T319 && T318;
  assign T318 = lockPortHadReadyRequest || lockPort_req_valid;
  assign T319 = ! AllOffloadsReady;
  assign T320 = lockPort_req_ready || lock_ready_received;
  assign T321 = T323 && T322;
  assign T322 = lock_ready_received || lockPort_req_ready;
  assign lockPort_req_ready = mainOff_lock_req_ready;
  assign T323 = ! AllOffloadsReady;
  assign T324 = T331 || T325;
  assign T325 = T327 && T326;
  assign T326 = ! memPort_req_valid;
  assign T327 = ! memPortHadReadyRequest;
  assign T328 = T330 && T329;
  assign T329 = memPortHadReadyRequest || memPort_req_valid;
  assign T330 = ! AllOffloadsReady;
  assign T331 = memPort_req_ready || mem_ready_received;
  assign T332 = T334 && T333;
  assign T333 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign T334 = ! AllOffloadsReady;
  assign T335 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T336;
  assign T336 = T337[8'ha5/* 165*/:8'h86/* 134*/];
  assign T337 = T481 ? T476 : T338;
  assign T338 = {T475, T474, T473, T472, T339};
  assign T339 = T340[2'h3/* 3*/:1'h0/* 0*/];
  assign T340 = T468 ? T454 : T341;
  assign T341 = {T453, T452, T451, T450, T342};
  assign T342 = T343[2'h3/* 3*/:1'h0/* 0*/];
  assign T343 = T446 ? T441 : T344;
  assign T344 = {T440, T439, T438, T437, T345};
  assign T345 = T346[2'h3/* 3*/:1'h0/* 0*/];
  assign T346 = T433 ? T348 : T347;
  assign T347 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T348 = {memReq4_addr, memReq4_rw, memReq4_cached, memReq4_data, memReq4_size};
  assign memReq4_size = 4'h8/* 8*/;
  assign memReq4_data = T349;
  assign T349 = {64'h0/* 0*/, T350};
  assign T350 = T415 | T351;
  assign T351 = rank_1 & T352;
  assign T352 = {7'h40/* 64*/{T8}};
  assign T353 = T251 || T249;
  assign T354 = T249 ? T395 : T355;
  assign T355 = T251 ? T357 : T356;
  assign T356 = {64'h0/* 0*/, rank_1};
  assign T357 = T386 | T358;
  assign T358 = memRep_1_data & T359;
  assign T359 = {8'h80/* 128*/{T122}};
  assign T360 = T361 || T247;
  assign T361 = T362 || T251;
  assign T362 = T255 || T253;
  assign T363 = T383 ? T364 : memRep_1_data;
  assign T364 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T380 ? T379 : T365;
  assign T365 = {T366};
  assign T366 = T374 | T367;
  assign T367 = memPortReplyStorage_1_data & T368;
  assign T368 = {8'h80/* 128*/{T122}};
  assign T369 = memPort_rep_valid && T370;
  assign T370 = T371[1'h1/* 1*/];
  assign T371 = T372[1'h1/* 1*/:1'h0/* 0*/];
  assign T372 = 2'h1/* 1*/ << memPort_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T373 = T369 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign T374 = memPortReplyStorage_0_data & T375;
  assign T375 = {8'h80/* 128*/{T133}};
  assign T376 = memPort_rep_valid && T377;
  assign T377 = T371[1'h0/* 0*/];
  assign T378 = T376 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T379 = {memPort_rep_bits_data};
  assign T380 = memPort_rep_valid && T381;
  assign T381 = T382 == memPort_rep_tag;
  assign T382 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T383 = T384 || T247;
  assign T384 = T385 || T251;
  assign T385 = T255 || T253;
  assign T386 = memRep_0_data & T387;
  assign T387 = {8'h80/* 128*/{T133}};
  assign T388 = T389 || T143;
  assign T389 = T390 || T155;
  assign T390 = T167 || T161;
  assign T391 = T392 ? T364 : memRep_0_data;
  assign T392 = T393 || T143;
  assign T393 = T394 || T155;
  assign T394 = T167 || T161;
  assign T395 = {64'h0/* 0*/, addOut_out};
  assign addOut_out = T396;
  assign T396 = addPortReplyValue[6'h3f/* 63*/:1'h0/* 0*/];
  assign addPortReplyValue = T412 ? T411 : T397;
  assign T397 = {T398};
  assign T398 = T406 | T399;
  assign T399 = addPortReplyStorage_1_out & T400;
  assign T400 = {7'h40/* 64*/{T122}};
  assign T401 = addPort_rep_valid && T402;
  assign T402 = T403[1'h1/* 1*/];
  assign T403 = T404[1'h1/* 1*/:1'h0/* 0*/];
  assign T404 = 2'h1/* 1*/ << addPort_rep_tag;
  assign T405 = T401 ? addPort_rep_bits_out : addPortReplyStorage_1_out;
  assign addPort_rep_bits_out = mainOff_add_rep_bits_out;
  assign T406 = addPortReplyStorage_0_out & T407;
  assign T407 = {7'h40/* 64*/{T133}};
  assign T408 = addPort_rep_valid && T409;
  assign T409 = T403[1'h0/* 0*/];
  assign T410 = T408 ? addPort_rep_bits_out : addPortReplyStorage_0_out;
  assign T411 = {addPort_rep_bits_out};
  assign T412 = addPort_rep_valid && T413;
  assign T413 = T414 == addPort_rep_tag;
  assign T414 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T415 = rank_0 & T416;
  assign T416 = {7'h40/* 64*/{T41}};
  assign T417 = T155 || T149;
  assign T418 = T149 ? T421 : T419;
  assign T419 = T155 ? T357 : T420;
  assign T420 = {64'h0/* 0*/, rank_0};
  assign T421 = {64'h0/* 0*/, addOut_out};
  assign memReq4_rw = 1'h1/* 1*/;
  assign memReq4_addr = T422;
  assign T422 = T423[5'h1f/* 31*/:1'h0/* 0*/];
  assign T423 = 56'h1000000/* 16777216*/ + T424;
  assign T424 = {21'h0/* 0*/, T425};
  assign T425 = T426 << 32'h3/* 3*/;
  assign T426 = T430 | T427;
  assign T427 = inputReg_1_pageId & T428;
  assign T428 = {6'h20/* 32*/{T8}};
  assign T429 = T184 ? io_in_bits_pageId : inputReg_1_pageId;
  assign T430 = inputReg_0_pageId & T431;
  assign T431 = {6'h20/* 32*/{T41}};
  assign T432 = T192 ? io_in_bits_pageId : inputReg_0_pageId;
  assign T433 = T436 && T434;
  assign T434 = T5 == T435;
  assign T435 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T436 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T437 = T346[8'h83/* 131*/:3'h4/* 4*/];
  assign T438 = T346[8'h84/* 132*/];
  assign T439 = T346[8'h85/* 133*/];
  assign T440 = T346[8'ha5/* 165*/:8'h86/* 134*/];
  assign T441 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h8/* 8*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T442;
  assign T442 = T443[5'h1f/* 31*/:1'h0/* 0*/];
  assign T443 = 56'h1000000/* 16777216*/ + T444;
  assign T444 = {21'h0/* 0*/, T445};
  assign T445 = T426 << 32'h3/* 3*/;
  assign T446 = T449 && T447;
  assign T447 = T5 == T448;
  assign T448 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T449 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T450 = T343[8'h83/* 131*/:3'h4/* 4*/];
  assign T451 = T343[8'h84/* 132*/];
  assign T452 = T343[8'h85/* 133*/];
  assign T453 = T343[8'ha5/* 165*/:8'h86/* 134*/];
  assign T454 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h4/* 4*/;
  assign memReq2_data = T455;
  assign T455 = T459 ^ T456;
  assign T456 = {96'h0/* 0*/, T457};
  assign T457 = 32'h1/* 1*/ << T458;
  assign T458 = T426 & 32'h1f/* 31*/;
  assign T459 = T462 | T460;
  assign T460 = memRep_1_data & T461;
  assign T461 = {8'h80/* 128*/{T8}};
  assign T462 = memRep_0_data & T463;
  assign T463 = {8'h80/* 128*/{T41}};
  assign memReq2_rw = 1'h1/* 1*/;
  assign memReq2_addr = T464;
  assign T464 = T465[5'h1f/* 31*/:1'h0/* 0*/];
  assign T465 = 59'h8000000/* 134217728*/ + T466;
  assign T466 = {27'h0/* 0*/, T467};
  assign T467 = T426 >> 32'h3/* 3*/;
  assign T468 = T471 && T469;
  assign T469 = T5 == T470;
  assign T470 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T471 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T472 = T340[8'h83/* 131*/:3'h4/* 4*/];
  assign T473 = T340[8'h84/* 132*/];
  assign T474 = T340[8'h85/* 133*/];
  assign T475 = T340[8'ha5/* 165*/:8'h86/* 134*/];
  assign T476 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h4/* 4*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T477;
  assign T477 = T478[5'h1f/* 31*/:1'h0/* 0*/];
  assign T478 = 59'h8000000/* 134217728*/ + T479;
  assign T479 = {27'h0/* 0*/, T480};
  assign T480 = T426 >> 32'h3/* 3*/;
  assign T481 = T484 && T482;
  assign T482 = T5 == T483;
  assign T483 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T484 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T485;
  assign T485 = T337[2'h3/* 3*/:1'h0/* 0*/];
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T486;
  assign T486 = T337[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T487;
  assign T487 = T337[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T488;
  assign T488 = T337[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T489;
  assign T489 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T490 = ! T491;
  assign T491 = T492 == 5'h1/* 1*/;
  assign T492 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T493 = mem_valid_received_0 & T41;
  assign T494 = T499 && T495;
  assign T495 = mem_valid_received_0 || T496;
  assign T496 = memPort_rep_valid && T497;
  assign T497 = memPort_rep_tag == T498;
  assign T498 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T499 = ! T500;
  assign T500 = T501 == 5'h0/* 0*/;
  assign T501 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T502 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T503 = 5'h1/* 1*/ == T504;
  assign T504 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T505 = ! T506;
  assign T506 = T507 == 5'h1/* 1*/;
  assign T507 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T508 = T509 || mem_valid_received_1;
  assign T509 = memPort_rep_valid && T510;
  assign T510 = memPort_rep_tag == T511;
  assign T511 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T512 = subStateTh_1 == 1'h1/* 1*/;
  assign T513 = T566 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T514;
  assign T514 = T529 && T515;
  assign T515 = T525 || T516;
  assign T516 = ! addPortHadValidRequest_0;
  assign T517 = T522 && T518;
  assign T518 = addPortHadValidRequest_0 || T519;
  assign T519 = T520 && addPort_req_valid;
  assign T520 = 5'h0/* 0*/ == T521;
  assign T521 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T522 = ! T523;
  assign T523 = T524 == 5'h0/* 0*/;
  assign T524 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T525 = T526 || add_valid_received_0;
  assign T526 = addPort_rep_valid && T527;
  assign T527 = addPort_rep_tag == T528;
  assign T528 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T529 = T552 && T530;
  assign T530 = T540 || T531;
  assign T531 = ! lockPortHadValidRequest_0;
  assign T532 = T537 && T533;
  assign T533 = lockPortHadValidRequest_0 || T534;
  assign T534 = T535 && lockPort_req_valid;
  assign T535 = 5'h0/* 0*/ == T536;
  assign T536 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T537 = ! T538;
  assign T538 = T539 == 5'h0/* 0*/;
  assign T539 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T540 = T549 || lock_valid_received_0;
  assign T541 = T546 && T542;
  assign T542 = lock_valid_received_0 || T543;
  assign T543 = lockPort_rep_valid && T544;
  assign T544 = lockPort_rep_tag == T545;
  assign T545 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T546 = ! T547;
  assign T547 = T548 == 5'h0/* 0*/;
  assign T548 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T549 = lockPort_rep_valid && T550;
  assign T550 = lockPort_rep_tag == T551;
  assign T551 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T552 = T562 || T553;
  assign T553 = ! memPortHadValidRequest_0;
  assign T554 = T559 && T555;
  assign T555 = memPortHadValidRequest_0 || T556;
  assign T556 = T557 && memPort_req_valid;
  assign T557 = 5'h0/* 0*/ == T558;
  assign T558 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T559 = ! T560;
  assign T560 = T561 == 5'h0/* 0*/;
  assign T561 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T562 = T563 || mem_valid_received_0;
  assign T563 = memPort_rep_valid && T564;
  assign T564 = memPort_rep_tag == T565;
  assign T565 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T566 = subStateTh_0 == 1'h1/* 1*/;
  assign T567 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T568 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T569 = T571 && T570;
  assign T570 = State_1 != 8'hff/* 255*/;
  assign T571 = T573 && T572;
  assign T572 = State_1 != 8'h0/* 0*/;
  assign T573 = AllOffloadsReady && T574;
  assign T574 = T575 == rThreadEncoder_io_chosen;
  assign T575 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T576 = subStateTh_0 == 1'h0/* 0*/;
  assign T577 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T578 = State_0 & T579;
  assign T579 = {4'h8/* 8*/{T41}};
  assign T580 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T581 = T584 && T582;
  assign T582 = T5 == T583;
  assign T583 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T584 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T585 = T590 && T586;
  assign T586 = ! T587;
  assign T587 = T589 | T588;
  assign T588 = lock_valid_received_1 & T8;
  assign T589 = lock_valid_received_0 & T41;
  assign T590 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_lock_req_tag = lockPort_req_tag;
  assign lockPort_req_tag = T591;
  assign T591 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign io_out_tag = T592;
  assign T592 = T596 | T593;
  assign T593 = inputTag_1 & T594;
  assign T594 = {4'ha/* 10*/{T8}};
  assign T595 = T184 ? io_in_tag : inputTag_1;
  assign T596 = inputTag_0 & T597;
  assign T597 = {4'ha/* 10*/{T41}};
  assign T598 = T192 ? io_in_tag : inputTag_0;
  RREncode_50 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T576 ),
       .io_valid_1( T11 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T577 ));
  RREncode_51 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T513 ),
       .io_valid_1( T15 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T567 ));
  RREncode_52 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T286 ),
       .io_valid_1( T118 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T335 ));

  always @(posedge clk) begin
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T12;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T19;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T31;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T42;
    lockPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T63;
    lock_valid_received_1 <= reset ? 1'h0/* 0*/ : T72;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T85;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T112;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T120) begin
      State_1 <= T264;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T134) begin
      State_0 <= T211;
    end
    if(T184) begin
      inputReg_1_done <= T190;
    end
    if(T192) begin
      inputReg_0_done <= T194;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      EmitReturnState_1 <= T228;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T232) begin
      EmitReturnState_0 <= T233;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T289;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T305;
    add_ready_received <= reset ? 1'h0/* 0*/ : T309;
    lockPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T317;
    lock_ready_received <= reset ? 1'h0/* 0*/ : T321;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T328;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T332;
    if(T353) begin
      rank_1 <= T354;
    end
    if(T360) begin
      memRep_1_data <= T363;
    end
    if(T369) begin
      memPortReplyStorage_1_data <= T373;
    end
    if(T376) begin
      memPortReplyStorage_0_data <= T378;
    end
    if(T388) begin
      memRep_0_data <= T391;
    end
    if(T401) begin
      addPortReplyStorage_1_out <= T405;
    end
    if(T408) begin
      addPortReplyStorage_0_out <= T410;
    end
    if(T417) begin
      rank_0 <= T418;
    end
    if(T184) begin
      inputReg_1_pageId <= T429;
    end
    if(T192) begin
      inputReg_0_pageId <= T432;
    end
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T494;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T517;
    lockPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T532;
    lock_valid_received_0 <= reset ? 1'h0/* 0*/ : T541;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T554;
    if(T184) begin
      inputTag_1 <= T595;
    end
    if(T192) begin
      inputTag_0 <= T598;
    end
  end
endmodule

module gPipe_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_7 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_19(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag,
    input  io_off_lock_req_ready,
    output io_off_lock_req_valid,
    output[31:0] io_off_lock_req_bits_id,
    output io_off_lock_req_bits_op,
    output[9:0] io_off_lock_req_tag,
    output io_off_lock_rep_ready,
    input  io_off_lock_rep_valid,
    input  io_off_lock_rep_bits_out,
    input [9:0] io_off_lock_rep_tag);

  wire mainComp_mainOff_lock_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire mainComp_mainOff_mem_req_valid;
  wire mainComp_mainOff_lock_rep_ready;
  wire mainComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_mainOff_lock_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_off_lock_req_valid = mainComp_mainOff_lock_req_valid;
  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_off_lock_rep_ready = mainComp_mainOff_lock_rep_ready;
  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_off_lock_req_tag = mainComp_mainOff_lock_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateWriter_2 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_lock_req_ready( io_off_lock_req_ready ),
       .mainOff_lock_req_valid( mainComp_mainOff_lock_req_valid ),
       .mainOff_lock_req_bits_id(  ),
       .mainOff_lock_req_bits_op(  ),
       .mainOff_lock_req_tag( mainComp_mainOff_lock_req_tag ),
       .mainOff_lock_rep_ready( mainComp_mainOff_lock_rep_ready ),
       .mainOff_lock_rep_valid( io_off_lock_rep_valid ),
       .mainOff_lock_rep_bits_out(  ),
       .mainOff_lock_rep_tag( io_off_lock_rep_tag ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_6 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_53(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_54(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module RREncode_55(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg[0:0] last_grant;
  wire T7;
  wire outValid;
  wire[1:0] T8;
  wire[1:0] T9;

  assign io_chosen = choose;
  assign choose = T5 ? T4 : T0;
  assign T0 = io_valid_0 ? T3 : T1;
  assign T1 = io_valid_1 ? T2 : 2'h2/* 2*/;
  assign T2 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T3 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = io_valid_1 && T6;
  assign T6 = 1'h1/* 1*/ > last_grant;
  assign T7 = outValid && io_ready;
  assign outValid = io_valid_0 || io_valid_1;
  assign T8 = T7 ? choose : T9;
  assign T9 = {1'h0/* 0*/, last_grant};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0/* 0*/;
    end else if(T7) begin
      last_grant <= T8;
    end
  end
endmodule

module updateWriter_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_lock_req_ready,
    output mainOff_lock_req_valid,
    output[31:0] mainOff_lock_req_bits_id,
    output mainOff_lock_req_bits_op,
    output[9:0] mainOff_lock_req_tag,
    output mainOff_lock_rep_ready,
    input  mainOff_lock_rep_valid,
    input  mainOff_lock_rep_bits_out,
    input [9:0] mainOff_lock_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_1;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[4:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_1;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_1;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[4:0] T24;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_1;
  wire T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire AllOffloadsReady;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg[0:0] addPortHadReadyRequest;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg[0:0] add_ready_received;
  wire T46;
  wire T47;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire lockPort_req_valid;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[7:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  reg[0:0] lock_valid_received_1;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[9:0] T71;
  wire[9:0] lockPort_rep_tag;
  wire lockPort_rep_ready;
  wire memPort_req_valid;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[7:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[7:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[7:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire[7:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg[0:0] mem_valid_received_1;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[9:0] T100;
  wire[9:0] memPort_rep_tag;
  wire memPort_rep_valid;
  wire T101;
  wire T102;
  wire[4:0] T103;
  wire T104;
  wire T105;
  reg[0:0] mem_valid_received_0;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[9:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[3:0] memPort_req_bits_size;
  wire[3:0] T118;
  wire[165:0] T119;
  wire[165:0] T120;
  wire[3:0] T121;
  wire[165:0] T122;
  wire[165:0] T123;
  wire[3:0] T124;
  wire[165:0] T125;
  wire[165:0] T126;
  wire[3:0] T127;
  wire[165:0] T128;
  wire[165:0] T129;
  wire[165:0] T130;
  wire[3:0] memReq4_size;
  wire[127:0] memReq4_data;
  wire[127:0] T131;
  wire[63:0] T132;
  wire[63:0] T133;
  wire[63:0] T134;
  reg[63:0] rank_1;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[7:0] T139;
  wire[7:0] T140;
  wire[7:0] T141;
  wire[7:0] T142;
  wire[7:0] T143;
  wire[7:0] T144;
  wire T145;
  reg[7:0] State_0;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[7:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire[7:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[7:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire[7:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[7:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire[7:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  reg[0:0] inputReg_1_done;
  wire T196;
  wire T197;
  wire[1:0] T198;
  wire[4:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  reg[0:0] inputReg_0_done;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire[7:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[7:0] T220;
  wire[7:0] T221;
  wire[7:0] T222;
  wire[7:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  wire[7:0] T226;
  wire[7:0] T227;
  wire[7:0] T228;
  wire[7:0] T229;
  wire[7:0] T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  reg[7:0] EmitReturnState_1;
  wire T235;
  wire T236;
  wire[7:0] T237;
  wire T238;
  wire[7:0] T239;
  wire[7:0] T240;
  reg[7:0] EmitReturnState_0;
  wire T241;
  wire[7:0] T242;
  wire T243;
  wire[7:0] T244;
  wire[7:0] T245;
  wire[7:0] T246;
  wire[7:0] T247;
  wire[7:0] T248;
  wire[7:0] T249;
  wire[7:0] T250;
  wire[7:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire[127:0] T255;
  wire[127:0] T256;
  wire[127:0] T257;
  wire[127:0] T258;
  wire[127:0] T259;
  wire[127:0] T260;
  reg[127:0] memRep_1_data;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire[127:0] T267;
  wire[127:0] T268;
  wire[127:0] memPortReplyValue;
  wire[127:0] T269;
  wire[127:0] T270;
  wire[127:0] T271;
  wire[127:0] T272;
  reg[127:0] memPortReplyStorage_1_data;
  wire T273;
  wire T274;
  wire[1:0] T275;
  wire[1024:0] T276;
  wire[127:0] T277;
  wire[127:0] memPort_rep_bits_data;
  wire[31:0] memPort_req_bits_addr;
  wire[31:0] T278;
  wire[127:0] T279;
  wire[127:0] T280;
  reg[127:0] memPortReplyStorage_0_data;
  wire T281;
  wire T282;
  wire[127:0] T283;
  wire[127:0] T284;
  wire T285;
  wire T286;
  wire[9:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[127:0] T291;
  wire[127:0] T292;
  reg[127:0] memRep_0_data;
  wire T293;
  wire T294;
  wire T295;
  wire[127:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire[127:0] T300;
  wire[63:0] addOut_out;
  wire[63:0] T301;
  wire[63:0] addPortReplyValue;
  wire[63:0] T302;
  wire[63:0] T303;
  wire[63:0] T304;
  wire[63:0] T305;
  reg[63:0] addPortReplyStorage_1_out;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire[1024:0] T309;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T310;
  wire addPort_rep_valid;
  wire[63:0] T311;
  wire[63:0] addPort_rep_bits_out;
  wire[63:0] T312;
  wire[63:0] T313;
  reg[63:0] addPortReplyStorage_0_out;
  wire T314;
  wire T315;
  wire[63:0] T316;
  wire[63:0] T317;
  wire T318;
  wire T319;
  wire[9:0] T320;
  wire[63:0] T321;
  wire[63:0] T322;
  reg[63:0] rank_0;
  wire T323;
  wire[127:0] T324;
  wire[127:0] T325;
  wire[127:0] T326;
  wire[127:0] T327;
  wire memReq4_cached;
  wire memReq4_rw;
  wire[31:0] memReq4_addr;
  wire[31:0] T328;
  wire[55:0] T329;
  wire[55:0] T330;
  wire[34:0] T331;
  wire[31:0] T332;
  wire[31:0] T333;
  wire[31:0] T334;
  reg[31:0] inputReg_1_pageId;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  reg[31:0] inputReg_0_pageId;
  wire[31:0] T338;
  wire T339;
  wire T340;
  wire[7:0] T341;
  wire T342;
  wire[127:0] T343;
  wire T344;
  wire T345;
  wire[31:0] T346;
  wire[165:0] T347;
  wire[3:0] memReq3_size;
  wire[127:0] memReq3_data;
  wire memReq3_cached;
  wire memReq3_rw;
  wire[31:0] memReq3_addr;
  wire[31:0] T348;
  wire[55:0] T349;
  wire[55:0] T350;
  wire[34:0] T351;
  wire T352;
  wire T353;
  wire[7:0] T354;
  wire T355;
  wire[127:0] T356;
  wire T357;
  wire T358;
  wire[31:0] T359;
  wire[165:0] T360;
  wire[3:0] memReq2_size;
  wire[127:0] memReq2_data;
  wire[127:0] T361;
  wire[127:0] T362;
  wire[31:0] T363;
  wire[31:0] T364;
  wire[127:0] T365;
  wire[127:0] T366;
  wire[127:0] T367;
  wire[127:0] T368;
  wire[127:0] T369;
  wire memReq2_cached;
  wire memReq2_rw;
  wire[31:0] memReq2_addr;
  wire[31:0] T370;
  wire[58:0] T371;
  wire[58:0] T372;
  wire[31:0] T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire[127:0] T378;
  wire T379;
  wire T380;
  wire[31:0] T381;
  wire[165:0] T382;
  wire[3:0] memReq1_size;
  wire[127:0] memReq1_data;
  wire memReq1_cached;
  wire memReq1_rw;
  wire[31:0] memReq1_addr;
  wire[31:0] T383;
  wire[58:0] T384;
  wire[58:0] T385;
  wire[31:0] T386;
  wire T387;
  wire T388;
  wire[7:0] T389;
  wire T390;
  wire[127:0] memPort_req_bits_data;
  wire[127:0] T391;
  wire memPort_req_bits_cached;
  wire T392;
  wire memPort_req_bits_rw;
  wire T393;
  wire memPort_rep_ready;
  wire[9:0] memPort_req_tag;
  wire[9:0] T394;
  wire[9:0] lockPort_req_tag;
  wire[9:0] T395;
  wire lockPort_rep_valid;
  wire T396;
  wire T397;
  wire[4:0] T398;
  wire T399;
  reg[0:0] lock_valid_received_0;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[9:0] T404;
  wire T405;
  wire T406;
  wire[4:0] T407;
  wire T408;
  wire T409;
  reg[0:0] lockPortHadReadyRequest;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  reg[0:0] lock_ready_received;
  wire T414;
  wire T415;
  wire lockPort_req_ready;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] memPortHadReadyRequest;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  reg[0:0] mem_ready_received;
  wire T425;
  wire T426;
  wire memPort_req_ready;
  wire T427;
  wire T428;
  reg[0:0] subStateTh_0;
  wire T429;
  wire T430;
  wire T431;
  wire[1:0] T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire[1:0] T439;
  wire T440;
  wire[7:0] T441;
  wire[7:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  reg[0:0] add_valid_received_1;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[9:0] T452;
  wire T453;
  wire T454;
  wire[4:0] T455;
  wire T456;
  reg[0:0] add_valid_received_0;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire[9:0] T461;
  wire T462;
  wire T463;
  wire[4:0] T464;
  wire T465;
  wire T466;
  wire[4:0] T467;
  wire T468;
  wire T469;
  wire[4:0] T470;
  wire T471;
  wire T472;
  wire T473;
  wire[9:0] T474;
  wire T475;
  wire T476;
  wire T477;
  reg[0:0] lockPortHadValidRequest_1;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire[4:0] T482;
  wire T483;
  wire T484;
  wire[4:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[9:0] T489;
  wire T490;
  wire T491;
  reg[0:0] memPortHadValidRequest_1;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire[4:0] T496;
  wire T497;
  wire T498;
  wire[4:0] T499;
  wire T500;
  wire T501;
  wire T502;
  wire[9:0] T503;
  wire T504;
  wire T505;
  wire AllOffloadsValid_0;
  wire T506;
  wire T507;
  wire T508;
  reg[0:0] addPortHadValidRequest_0;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire[4:0] T513;
  wire T514;
  wire T515;
  wire[4:0] T516;
  wire T517;
  wire T518;
  wire T519;
  wire[9:0] T520;
  wire T521;
  wire T522;
  wire T523;
  reg[0:0] lockPortHadValidRequest_0;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire[4:0] T528;
  wire T529;
  wire T530;
  wire[4:0] T531;
  wire T532;
  wire T533;
  wire T534;
  wire[9:0] T535;
  wire T536;
  wire T537;
  reg[0:0] memPortHadValidRequest_0;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[4:0] T542;
  wire T543;
  wire T544;
  wire[4:0] T545;
  wire T546;
  wire T547;
  wire T548;
  wire[9:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire[7:0] T570;
  wire[7:0] T571;
  wire[7:0] T572;
  wire[7:0] T573;
  wire[7:0] T574;
  wire[7:0] T575;
  wire[7:0] T576;
  wire[7:0] T577;
  wire[7:0] T578;
  wire[7:0] T579;
  wire[7:0] T580;
  wire[7:0] T581;
  wire[7:0] T582;
  wire[7:0] T583;
  wire[7:0] T584;
  wire[7:0] T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[9:0] T592;
  wire[9:0] T593;
  wire[9:0] T594;
  reg[9:0] inputTag_1;
  wire[9:0] T595;
  wire[9:0] T596;
  wire[9:0] T597;
  reg[9:0] inputTag_0;
  wire[9:0] T598;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T1 = T587 && T2;
  assign T2 = State_1 == 8'h0/* 0*/;
  assign T3 = T552 || T4;
  assign T4 = T148 && T5;
  assign T5 = T6[1'h1/* 1*/];
  assign T6 = T7[1'h1/* 1*/:1'h0/* 0*/];
  assign T7 = 2'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T504 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T9;
  assign T9 = T475 && T10;
  assign T10 = T471 || T11;
  assign T11 = ! addPortHadValidRequest_1;
  assign T12 = T468 && T13;
  assign T13 = addPortHadValidRequest_1 || T14;
  assign T14 = T466 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T444 && T16;
  assign T16 = T443 && T17;
  assign T17 = T19 == T18;
  assign T18 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T19 = T441 | T20;
  assign T20 = State_1 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23[1'h1/* 1*/];
  assign T23 = T24[1'h1/* 1*/:1'h0/* 0*/];
  assign T24 = 2'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_1 == 1'h0/* 0*/;
  assign T26 = T30 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_1;
  assign T28 = T29 == vThreadEncoder_io_chosen;
  assign T29 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T30 = T32 && T31;
  assign T31 = State_1 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_1 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = T36 == rThreadEncoder_io_chosen;
  assign T36 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign AllOffloadsReady = T37;
  assign T37 = T49 && T38;
  assign T38 = T45 || T39;
  assign T39 = T41 && T40;
  assign T40 = ! addPort_req_valid;
  assign T41 = ! addPortHadReadyRequest;
  assign T42 = T44 && T43;
  assign T43 = addPortHadReadyRequest || addPort_req_valid;
  assign T44 = ! AllOffloadsReady;
  assign T45 = addPort_req_ready || add_ready_received;
  assign T46 = T48 && T47;
  assign T47 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T48 = ! AllOffloadsReady;
  assign T49 = T417 && T50;
  assign T50 = T413 || T51;
  assign T51 = T409 && T52;
  assign T52 = ! lockPort_req_valid;
  assign lockPort_req_valid = T53;
  assign T53 = T63 && T54;
  assign T54 = T59 || T55;
  assign T55 = T58 && T56;
  assign T56 = T19 == T57;
  assign T57 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T58 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T59 = T62 && T60;
  assign T60 = T19 == T61;
  assign T61 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T63 = T408 && T64;
  assign T64 = ! T65;
  assign T65 = T399 | T66;
  assign T66 = lock_valid_received_1 & T22;
  assign T67 = T396 && T68;
  assign T68 = lock_valid_received_1 || T69;
  assign T69 = lockPort_rep_valid && T70;
  assign T70 = lockPort_rep_tag == T71;
  assign T71 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign lockPort_rep_tag = mainOff_lock_rep_tag;
  assign mainOff_lock_req_valid = lockPort_req_valid;
  assign mainOff_lock_rep_ready = lockPort_rep_ready;
  assign lockPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_valid = memPort_req_valid;
  assign memPort_req_valid = T72;
  assign T72 = T92 && T73;
  assign T73 = T78 || T74;
  assign T74 = T77 && T75;
  assign T75 = T19 == T76;
  assign T76 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T77 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T78 = T83 || T79;
  assign T79 = T82 && T80;
  assign T80 = T19 == T81;
  assign T81 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T82 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T83 = T88 || T84;
  assign T84 = T87 && T85;
  assign T85 = T19 == T86;
  assign T86 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T87 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T88 = T91 && T89;
  assign T89 = T19 == T90;
  assign T90 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T91 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T92 = T114 && T93;
  assign T93 = ! T94;
  assign T94 = T104 | T95;
  assign T95 = mem_valid_received_1 & T22;
  assign T96 = T101 && T97;
  assign T97 = mem_valid_received_1 || T98;
  assign T98 = memPort_rep_valid && T99;
  assign T99 = memPort_rep_tag == T100;
  assign T100 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign memPort_rep_tag = mainOff_mem_rep_tag;
  assign memPort_rep_valid = mainOff_mem_rep_valid;
  assign T101 = ! T102;
  assign T102 = T103 == 5'h1/* 1*/;
  assign T103 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T104 = mem_valid_received_0 & T105;
  assign T105 = T23[1'h0/* 0*/];
  assign T106 = T111 && T107;
  assign T107 = mem_valid_received_0 || T108;
  assign T108 = memPort_rep_valid && T109;
  assign T109 = memPort_rep_tag == T110;
  assign T110 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_valid = T115;
  assign T115 = T117 && T116;
  assign T116 = T19 == 8'hff/* 255*/;
  assign T117 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_size = memPort_req_bits_size;
  assign memPort_req_bits_size = T118;
  assign T118 = T119[2'h3/* 3*/:1'h0/* 0*/];
  assign T119 = T387 ? T382 : T120;
  assign T120 = {T381, T380, T379, T378, T121};
  assign T121 = T122[2'h3/* 3*/:1'h0/* 0*/];
  assign T122 = T374 ? T360 : T123;
  assign T123 = {T359, T358, T357, T356, T124};
  assign T124 = T125[2'h3/* 3*/:1'h0/* 0*/];
  assign T125 = T352 ? T347 : T126;
  assign T126 = {T346, T345, T344, T343, T127};
  assign T127 = T128[2'h3/* 3*/:1'h0/* 0*/];
  assign T128 = T339 ? T130 : T129;
  assign T129 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T130 = {memReq4_addr, memReq4_rw, memReq4_cached, memReq4_data, memReq4_size};
  assign memReq4_size = 4'h8/* 8*/;
  assign memReq4_data = T131;
  assign T131 = {64'h0/* 0*/, T132};
  assign T132 = T321 | T133;
  assign T133 = rank_1 & T134;
  assign T134 = {7'h40/* 64*/{T22}};
  assign T135 = T254 || T136;
  assign T136 = T137 && T5;
  assign T137 = T253 && T138;
  assign T138 = T140 == T139;
  assign T139 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T140 = T143 | T141;
  assign T141 = State_1 & T142;
  assign T142 = {4'h8/* 8*/{T5}};
  assign T143 = State_0 & T144;
  assign T144 = {4'h8/* 8*/{T145}};
  assign T145 = T6[1'h0/* 0*/];
  assign T146 = T152 || T147;
  assign T147 = T148 && T145;
  assign T148 = T151 && T149;
  assign T149 = T140 == T150;
  assign T150 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T151 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T152 = T158 || T153;
  assign T153 = T154 && T145;
  assign T154 = T157 && T155;
  assign T155 = T140 == T156;
  assign T156 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T157 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T158 = T164 || T159;
  assign T159 = T160 && T145;
  assign T160 = T163 && T161;
  assign T161 = T140 == T162;
  assign T162 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T163 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T164 = T166 || T165;
  assign T165 = T137 && T145;
  assign T166 = T172 || T167;
  assign T167 = T168 && T145;
  assign T168 = T171 && T169;
  assign T169 = T140 == T170;
  assign T170 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T171 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T172 = T178 || T173;
  assign T173 = T174 && T145;
  assign T174 = T177 && T175;
  assign T175 = T140 == T176;
  assign T176 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T177 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T178 = T184 || T179;
  assign T179 = T180 && T145;
  assign T180 = T183 && T181;
  assign T181 = T140 == T182;
  assign T182 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T183 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T184 = T190 || T185;
  assign T185 = T186 && T145;
  assign T186 = T189 && T187;
  assign T187 = T140 == T188;
  assign T188 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T189 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T190 = T211 || T191;
  assign T191 = T192 && T145;
  assign T192 = T207 && T193;
  assign T193 = ! T194;
  assign T194 = T203 | T195;
  assign T195 = inputReg_1_done & T5;
  assign T196 = T200 && T197;
  assign T197 = T198[1'h1/* 1*/];
  assign T198 = T199[1'h1/* 1*/:1'h0/* 0*/];
  assign T199 = 2'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T200 = T201 && io_in_valid;
  assign T201 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T202 = T196 ? io_in_bits_done : inputReg_1_done;
  assign T203 = inputReg_0_done & T145;
  assign T204 = T200 && T205;
  assign T205 = T198[1'h0/* 0*/];
  assign T206 = T204 ? io_in_bits_done : inputReg_0_done;
  assign T207 = T210 && T208;
  assign T208 = T140 == T209;
  assign T209 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T210 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T211 = T214 || T212;
  assign T212 = T213 && T145;
  assign T213 = T207 && T194;
  assign T214 = T204 || T215;
  assign T215 = T216 && T105;
  assign T216 = T217 && io_out_ready;
  assign T217 = T219 && T218;
  assign T218 = T19 == 8'hff/* 255*/;
  assign T219 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T220 = T252 ? 8'hff/* 255*/ : T221;
  assign T221 = T159 ? T251 : T222;
  assign T222 = T165 ? T250 : T223;
  assign T223 = T167 ? T249 : T224;
  assign T224 = T173 ? T248 : T225;
  assign T225 = T179 ? T247 : T226;
  assign T226 = T185 ? T246 : T227;
  assign T227 = T191 ? T245 : T228;
  assign T228 = T212 ? T244 : T229;
  assign T229 = T215 ? T232 : T230;
  assign T230 = T204 ? T231 : State_0;
  assign T231 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T232 = T239 | T233;
  assign T233 = EmitReturnState_1 & T234;
  assign T234 = {4'h8/* 8*/{T22}};
  assign T235 = T236 || T4;
  assign T236 = T154 && T5;
  assign T237 = T238 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T238 = T236 || T4;
  assign T239 = EmitReturnState_0 & T240;
  assign T240 = {4'h8/* 8*/{T105}};
  assign T241 = T153 || T147;
  assign T242 = T243 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T243 = T153 || T147;
  assign T244 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T245 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T246 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T247 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T248 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T249 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T250 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T251 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T252 = T153 || T147;
  assign T253 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T254 = T168 && T5;
  assign T255 = T136 ? T300 : T256;
  assign T256 = T254 ? T258 : T257;
  assign T257 = {64'h0/* 0*/, rank_1};
  assign T258 = T291 | T259;
  assign T259 = memRep_1_data & T260;
  assign T260 = {8'h80/* 128*/{T5}};
  assign T261 = T263 || T262;
  assign T262 = T160 && T5;
  assign T263 = T264 || T254;
  assign T264 = T266 || T265;
  assign T265 = T174 && T5;
  assign T266 = T180 && T5;
  assign T267 = T288 ? T268 : memRep_1_data;
  assign T268 = memPortReplyValue[7'h7f/* 127*/:1'h0/* 0*/];
  assign memPortReplyValue = T285 ? T284 : T269;
  assign T269 = {T270};
  assign T270 = T279 | T271;
  assign T271 = memPortReplyStorage_1_data & T272;
  assign T272 = {8'h80/* 128*/{T5}};
  assign T273 = memPort_rep_valid && T274;
  assign T274 = T275[1'h1/* 1*/];
  assign T275 = T276[1'h1/* 1*/:1'h0/* 0*/];
  assign T276 = 2'h1/* 1*/ << memPort_rep_tag;
  assign T277 = T273 ? memPort_rep_bits_data : memPortReplyStorage_1_data;
  assign memPort_rep_bits_data = mainOff_mem_rep_bits_data;
  assign mainOff_mem_req_bits_addr = memPort_req_bits_addr;
  assign memPort_req_bits_addr = T278;
  assign T278 = T119[8'ha5/* 165*/:8'h86/* 134*/];
  assign T279 = memPortReplyStorage_0_data & T280;
  assign T280 = {8'h80/* 128*/{T145}};
  assign T281 = memPort_rep_valid && T282;
  assign T282 = T275[1'h0/* 0*/];
  assign T283 = T281 ? memPort_rep_bits_data : memPortReplyStorage_0_data;
  assign T284 = {memPort_rep_bits_data};
  assign T285 = memPort_rep_valid && T286;
  assign T286 = T287 == memPort_rep_tag;
  assign T287 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T288 = T289 || T262;
  assign T289 = T290 || T254;
  assign T290 = T266 || T265;
  assign T291 = memRep_0_data & T292;
  assign T292 = {8'h80/* 128*/{T145}};
  assign T293 = T294 || T159;
  assign T294 = T295 || T167;
  assign T295 = T179 || T173;
  assign T296 = T297 ? T268 : memRep_0_data;
  assign T297 = T298 || T159;
  assign T298 = T299 || T167;
  assign T299 = T179 || T173;
  assign T300 = {64'h0/* 0*/, addOut_out};
  assign addOut_out = T301;
  assign T301 = addPortReplyValue[6'h3f/* 63*/:1'h0/* 0*/];
  assign addPortReplyValue = T318 ? T317 : T302;
  assign T302 = {T303};
  assign T303 = T312 | T304;
  assign T304 = addPortReplyStorage_1_out & T305;
  assign T305 = {7'h40/* 64*/{T5}};
  assign T306 = addPort_rep_valid && T307;
  assign T307 = T308[1'h1/* 1*/];
  assign T308 = T309[1'h1/* 1*/:1'h0/* 0*/];
  assign T309 = 2'h1/* 1*/ << addPort_rep_tag;
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T310;
  assign T310 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T311 = T306 ? addPort_rep_bits_out : addPortReplyStorage_1_out;
  assign addPort_rep_bits_out = mainOff_add_rep_bits_out;
  assign T312 = addPortReplyStorage_0_out & T313;
  assign T313 = {7'h40/* 64*/{T145}};
  assign T314 = addPort_rep_valid && T315;
  assign T315 = T308[1'h0/* 0*/];
  assign T316 = T314 ? addPort_rep_bits_out : addPortReplyStorage_0_out;
  assign T317 = {addPort_rep_bits_out};
  assign T318 = addPort_rep_valid && T319;
  assign T319 = T320 == addPort_rep_tag;
  assign T320 = {8'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T321 = rank_0 & T322;
  assign T322 = {7'h40/* 64*/{T105}};
  assign T323 = T167 || T165;
  assign T324 = T165 ? T327 : T325;
  assign T325 = T167 ? T258 : T326;
  assign T326 = {64'h0/* 0*/, rank_0};
  assign T327 = {64'h0/* 0*/, addOut_out};
  assign memReq4_rw = 1'h1/* 1*/;
  assign memReq4_addr = T328;
  assign T328 = T329[5'h1f/* 31*/:1'h0/* 0*/];
  assign T329 = 56'h1000000/* 16777216*/ + T330;
  assign T330 = {21'h0/* 0*/, T331};
  assign T331 = T332 << 32'h3/* 3*/;
  assign T332 = T336 | T333;
  assign T333 = inputReg_1_pageId & T334;
  assign T334 = {6'h20/* 32*/{T22}};
  assign T335 = T196 ? io_in_bits_pageId : inputReg_1_pageId;
  assign T336 = inputReg_0_pageId & T337;
  assign T337 = {6'h20/* 32*/{T105}};
  assign T338 = T204 ? io_in_bits_pageId : inputReg_0_pageId;
  assign T339 = T342 && T340;
  assign T340 = T19 == T341;
  assign T341 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T342 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T343 = T128[8'h83/* 131*/:3'h4/* 4*/];
  assign T344 = T128[8'h84/* 132*/];
  assign T345 = T128[8'h85/* 133*/];
  assign T346 = T128[8'ha5/* 165*/:8'h86/* 134*/];
  assign T347 = {memReq3_addr, memReq3_rw, memReq3_cached, memReq3_data, memReq3_size};
  assign memReq3_size = 4'h8/* 8*/;
  assign memReq3_rw = 1'h0/* 0*/;
  assign memReq3_addr = T348;
  assign T348 = T349[5'h1f/* 31*/:1'h0/* 0*/];
  assign T349 = 56'h1000000/* 16777216*/ + T350;
  assign T350 = {21'h0/* 0*/, T351};
  assign T351 = T332 << 32'h3/* 3*/;
  assign T352 = T355 && T353;
  assign T353 = T19 == T354;
  assign T354 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T355 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T356 = T125[8'h83/* 131*/:3'h4/* 4*/];
  assign T357 = T125[8'h84/* 132*/];
  assign T358 = T125[8'h85/* 133*/];
  assign T359 = T125[8'ha5/* 165*/:8'h86/* 134*/];
  assign T360 = {memReq2_addr, memReq2_rw, memReq2_cached, memReq2_data, memReq2_size};
  assign memReq2_size = 4'h4/* 4*/;
  assign memReq2_data = T361;
  assign T361 = T365 ^ T362;
  assign T362 = {96'h0/* 0*/, T363};
  assign T363 = 32'h1/* 1*/ << T364;
  assign T364 = T332 & 32'h1f/* 31*/;
  assign T365 = T368 | T366;
  assign T366 = memRep_1_data & T367;
  assign T367 = {8'h80/* 128*/{T22}};
  assign T368 = memRep_0_data & T369;
  assign T369 = {8'h80/* 128*/{T105}};
  assign memReq2_rw = 1'h1/* 1*/;
  assign memReq2_addr = T370;
  assign T370 = T371[5'h1f/* 31*/:1'h0/* 0*/];
  assign T371 = 59'h8000000/* 134217728*/ + T372;
  assign T372 = {27'h0/* 0*/, T373};
  assign T373 = T332 >> 32'h3/* 3*/;
  assign T374 = T377 && T375;
  assign T375 = T19 == T376;
  assign T376 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T377 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T378 = T122[8'h83/* 131*/:3'h4/* 4*/];
  assign T379 = T122[8'h84/* 132*/];
  assign T380 = T122[8'h85/* 133*/];
  assign T381 = T122[8'ha5/* 165*/:8'h86/* 134*/];
  assign T382 = {memReq1_addr, memReq1_rw, memReq1_cached, memReq1_data, memReq1_size};
  assign memReq1_size = 4'h4/* 4*/;
  assign memReq1_rw = 1'h0/* 0*/;
  assign memReq1_addr = T383;
  assign T383 = T384[5'h1f/* 31*/:1'h0/* 0*/];
  assign T384 = 59'h8000000/* 134217728*/ + T385;
  assign T385 = {27'h0/* 0*/, T386};
  assign T386 = T332 >> 32'h3/* 3*/;
  assign T387 = T390 && T388;
  assign T388 = T19 == T389;
  assign T389 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T390 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign mainOff_mem_req_bits_data = memPort_req_bits_data;
  assign memPort_req_bits_data = T391;
  assign T391 = T119[8'h83/* 131*/:3'h4/* 4*/];
  assign mainOff_mem_req_bits_cached = memPort_req_bits_cached;
  assign memPort_req_bits_cached = T392;
  assign T392 = T119[8'h84/* 132*/];
  assign mainOff_mem_req_bits_rw = memPort_req_bits_rw;
  assign memPort_req_bits_rw = T393;
  assign T393 = T119[8'h85/* 133*/];
  assign mainOff_mem_rep_ready = memPort_rep_ready;
  assign memPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_mem_req_tag = memPort_req_tag;
  assign memPort_req_tag = T394;
  assign T394 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mainOff_lock_req_tag = lockPort_req_tag;
  assign lockPort_req_tag = T395;
  assign T395 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign lockPort_rep_valid = mainOff_lock_rep_valid;
  assign T396 = ! T397;
  assign T397 = T398 == 5'h1/* 1*/;
  assign T398 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T399 = lock_valid_received_0 & T105;
  assign T400 = T405 && T401;
  assign T401 = lock_valid_received_0 || T402;
  assign T402 = lockPort_rep_valid && T403;
  assign T403 = lockPort_rep_tag == T404;
  assign T404 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T405 = ! T406;
  assign T406 = T407 == 5'h0/* 0*/;
  assign T407 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T408 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T409 = ! lockPortHadReadyRequest;
  assign T410 = T412 && T411;
  assign T411 = lockPortHadReadyRequest || lockPort_req_valid;
  assign T412 = ! AllOffloadsReady;
  assign T413 = lockPort_req_ready || lock_ready_received;
  assign T414 = T416 && T415;
  assign T415 = lock_ready_received || lockPort_req_ready;
  assign lockPort_req_ready = mainOff_lock_req_ready;
  assign T416 = ! AllOffloadsReady;
  assign T417 = T424 || T418;
  assign T418 = T420 && T419;
  assign T419 = ! memPort_req_valid;
  assign T420 = ! memPortHadReadyRequest;
  assign T421 = T423 && T422;
  assign T422 = memPortHadReadyRequest || memPort_req_valid;
  assign T423 = ! AllOffloadsReady;
  assign T424 = memPort_req_ready || mem_ready_received;
  assign T425 = T427 && T426;
  assign T426 = mem_ready_received || memPort_req_ready;
  assign memPort_req_ready = mainOff_mem_req_ready;
  assign T427 = ! AllOffloadsReady;
  assign T428 = subStateTh_0 == 1'h0/* 0*/;
  assign T429 = T433 ? 1'h1/* 1*/ : T430;
  assign T430 = T431 ? 1'h0/* 0*/ : subStateTh_0;
  assign T431 = T432 == vThreadEncoder_io_chosen;
  assign T432 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T433 = T435 && T434;
  assign T434 = State_0 != 8'hff/* 255*/;
  assign T435 = T437 && T436;
  assign T436 = State_0 != 8'h0/* 0*/;
  assign T437 = AllOffloadsReady && T438;
  assign T438 = T439 == rThreadEncoder_io_chosen;
  assign T439 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T440 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T441 = State_0 & T442;
  assign T442 = {4'h8/* 8*/{T105}};
  assign T443 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T444 = T465 && T445;
  assign T445 = ! T446;
  assign T446 = T456 | T447;
  assign T447 = add_valid_received_1 & T22;
  assign T448 = T453 && T449;
  assign T449 = add_valid_received_1 || T450;
  assign T450 = addPort_rep_valid && T451;
  assign T451 = addPort_rep_tag == T452;
  assign T452 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T453 = ! T454;
  assign T454 = T455 == 5'h1/* 1*/;
  assign T455 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T456 = add_valid_received_0 & T105;
  assign T457 = T462 && T458;
  assign T458 = add_valid_received_0 || T459;
  assign T459 = addPort_rep_valid && T460;
  assign T460 = addPort_rep_tag == T461;
  assign T461 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T462 = ! T463;
  assign T463 = T464 == 5'h0/* 0*/;
  assign T464 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T465 = rThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T466 = 5'h1/* 1*/ == T467;
  assign T467 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T468 = ! T469;
  assign T469 = T470 == 5'h1/* 1*/;
  assign T470 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T471 = T472 || add_valid_received_1;
  assign T472 = addPort_rep_valid && T473;
  assign T473 = addPort_rep_tag == T474;
  assign T474 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T475 = T490 && T476;
  assign T476 = T486 || T477;
  assign T477 = ! lockPortHadValidRequest_1;
  assign T478 = T483 && T479;
  assign T479 = lockPortHadValidRequest_1 || T480;
  assign T480 = T481 && lockPort_req_valid;
  assign T481 = 5'h1/* 1*/ == T482;
  assign T482 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T483 = ! T484;
  assign T484 = T485 == 5'h1/* 1*/;
  assign T485 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T486 = T487 || lock_valid_received_1;
  assign T487 = lockPort_rep_valid && T488;
  assign T488 = lockPort_rep_tag == T489;
  assign T489 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T490 = T500 || T491;
  assign T491 = ! memPortHadValidRequest_1;
  assign T492 = T497 && T493;
  assign T493 = memPortHadValidRequest_1 || T494;
  assign T494 = T495 && memPort_req_valid;
  assign T495 = 5'h1/* 1*/ == T496;
  assign T496 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T497 = ! T498;
  assign T498 = T499 == 5'h1/* 1*/;
  assign T499 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T500 = T501 || mem_valid_received_1;
  assign T501 = memPort_rep_valid && T502;
  assign T502 = memPort_rep_tag == T503;
  assign T503 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T504 = subStateTh_1 == 1'h1/* 1*/;
  assign T505 = T550 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T506;
  assign T506 = T521 && T507;
  assign T507 = T517 || T508;
  assign T508 = ! addPortHadValidRequest_0;
  assign T509 = T514 && T510;
  assign T510 = addPortHadValidRequest_0 || T511;
  assign T511 = T512 && addPort_req_valid;
  assign T512 = 5'h0/* 0*/ == T513;
  assign T513 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T514 = ! T515;
  assign T515 = T516 == 5'h0/* 0*/;
  assign T516 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T517 = T518 || add_valid_received_0;
  assign T518 = addPort_rep_valid && T519;
  assign T519 = addPort_rep_tag == T520;
  assign T520 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T521 = T536 && T522;
  assign T522 = T532 || T523;
  assign T523 = ! lockPortHadValidRequest_0;
  assign T524 = T529 && T525;
  assign T525 = lockPortHadValidRequest_0 || T526;
  assign T526 = T527 && lockPort_req_valid;
  assign T527 = 5'h0/* 0*/ == T528;
  assign T528 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T529 = ! T530;
  assign T530 = T531 == 5'h0/* 0*/;
  assign T531 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T532 = T533 || lock_valid_received_0;
  assign T533 = lockPort_rep_valid && T534;
  assign T534 = lockPort_rep_tag == T535;
  assign T535 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T536 = T546 || T537;
  assign T537 = ! memPortHadValidRequest_0;
  assign T538 = T543 && T539;
  assign T539 = memPortHadValidRequest_0 || T540;
  assign T540 = T541 && memPort_req_valid;
  assign T541 = 5'h0/* 0*/ == T542;
  assign T542 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T543 = ! T544;
  assign T544 = T545 == 5'h0/* 0*/;
  assign T545 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T546 = T547 || mem_valid_received_0;
  assign T547 = memPort_rep_valid && T548;
  assign T548 = memPort_rep_tag == T549;
  assign T549 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T550 = subStateTh_0 == 1'h1/* 1*/;
  assign T551 = vThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign T552 = T553 || T236;
  assign T553 = T554 || T262;
  assign T554 = T555 || T136;
  assign T555 = T556 || T254;
  assign T556 = T557 || T265;
  assign T557 = T558 || T266;
  assign T558 = T560 || T559;
  assign T559 = T186 && T5;
  assign T560 = T562 || T561;
  assign T561 = T192 && T5;
  assign T562 = T564 || T563;
  assign T563 = T213 && T5;
  assign T564 = T196 || T565;
  assign T565 = T216 && T22;
  assign T566 = T586 ? 8'hff/* 255*/ : T567;
  assign T567 = T262 ? T585 : T568;
  assign T568 = T136 ? T584 : T569;
  assign T569 = T254 ? T583 : T570;
  assign T570 = T265 ? T582 : T571;
  assign T571 = T266 ? T581 : T572;
  assign T572 = T559 ? T580 : T573;
  assign T573 = T561 ? T579 : T574;
  assign T574 = T563 ? T578 : T575;
  assign T575 = T565 ? T232 : T576;
  assign T576 = T196 ? T577 : State_1;
  assign T577 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T578 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T579 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T580 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T581 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T582 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T583 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T584 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T585 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T586 = T236 || T4;
  assign T587 = subStateTh_1 == 1'h0/* 0*/;
  assign T588 = T590 && T589;
  assign T589 = State_0 == 8'h0/* 0*/;
  assign T590 = subStateTh_0 == 1'h0/* 0*/;
  assign T591 = sThreadEncoder_io_chosen != 2'h2/* 2*/;
  assign io_out_tag = T592;
  assign T592 = T596 | T593;
  assign T593 = inputTag_1 & T594;
  assign T594 = {4'ha/* 10*/{T22}};
  assign T595 = T196 ? io_in_tag : inputTag_1;
  assign T596 = inputTag_0 & T597;
  assign T597 = {4'ha/* 10*/{T105}};
  assign T598 = T204 ? io_in_tag : inputTag_0;
  RREncode_53 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T428 ),
       .io_valid_1( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T440 ));
  RREncode_54 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T505 ),
       .io_valid_1( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T551 ));
  RREncode_55 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T588 ),
       .io_valid_1( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T591 ));

  always @(posedge clk) begin
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_1 <= T566;
    end
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T26;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T42;
    add_ready_received <= reset ? 1'h0/* 0*/ : T46;
    lock_valid_received_1 <= reset ? 1'h0/* 0*/ : T67;
    mem_valid_received_1 <= reset ? 1'h0/* 0*/ : T96;
    mem_valid_received_0 <= reset ? 1'h0/* 0*/ : T106;
    if(T135) begin
      rank_1 <= T255;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T146) begin
      State_0 <= T220;
    end
    if(T196) begin
      inputReg_1_done <= T202;
    end
    if(T204) begin
      inputReg_0_done <= T206;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T235) begin
      EmitReturnState_1 <= T237;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      EmitReturnState_0 <= T242;
    end
    if(T261) begin
      memRep_1_data <= T267;
    end
    if(T273) begin
      memPortReplyStorage_1_data <= T277;
    end
    if(T281) begin
      memPortReplyStorage_0_data <= T283;
    end
    if(T293) begin
      memRep_0_data <= T296;
    end
    if(T306) begin
      addPortReplyStorage_1_out <= T311;
    end
    if(T314) begin
      addPortReplyStorage_0_out <= T316;
    end
    if(T323) begin
      rank_0 <= T324;
    end
    if(T196) begin
      inputReg_1_pageId <= T335;
    end
    if(T204) begin
      inputReg_0_pageId <= T338;
    end
    lock_valid_received_0 <= reset ? 1'h0/* 0*/ : T400;
    lockPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T410;
    lock_ready_received <= reset ? 1'h0/* 0*/ : T414;
    memPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T421;
    mem_ready_received <= reset ? 1'h0/* 0*/ : T425;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T429;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T448;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T457;
    lockPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T478;
    memPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T492;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T509;
    lockPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T524;
    memPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T538;
    if(T196) begin
      inputTag_1 <= T595;
    end
    if(T204) begin
      inputTag_0 <= T598;
    end
  end
endmodule

module gPipe_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_8 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_20(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output pcOutN_valid,
    output pcOutN_bits_request,
    output[15:0] pcOutN_bits_moduleId,
    output[7:0] pcOutN_bits_portId,
    output[19:0] pcOutN_bits_pcValue,
    output[3:0] pcOutN_bits_pcType,
    input  io_off_mem_req_ready,
    output io_off_mem_req_valid,
    output[31:0] io_off_mem_req_bits_addr,
    output io_off_mem_req_bits_rw,
    output io_off_mem_req_bits_cached,
    output[127:0] io_off_mem_req_bits_data,
    output[3:0] io_off_mem_req_bits_size,
    output[9:0] io_off_mem_req_tag,
    output io_off_mem_rep_ready,
    input  io_off_mem_rep_valid,
    input [127:0] io_off_mem_rep_bits_data,
    input [9:0] io_off_mem_rep_tag,
    input  io_off_lock_req_ready,
    output io_off_lock_req_valid,
    output[31:0] io_off_lock_req_bits_id,
    output io_off_lock_req_bits_op,
    output[9:0] io_off_lock_req_tag,
    output io_off_lock_rep_ready,
    input  io_off_lock_rep_valid,
    input  io_off_lock_rep_bits_out,
    input [9:0] io_off_lock_rep_tag);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_mainOff_lock_req_valid;
  wire mainComp_mainOff_lock_rep_ready;
  wire mainComp_mainOff_mem_req_valid;
  wire mainComp_io_out_valid;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_mainOff_lock_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_off_lock_req_valid = mainComp_mainOff_lock_req_valid;
  assign io_off_lock_rep_ready = mainComp_mainOff_lock_rep_ready;
  assign io_off_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_off_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign io_off_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign io_off_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign io_off_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign io_off_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign io_off_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign io_off_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_off_lock_req_tag = mainComp_mainOff_lock_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  updateWriter_3 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( io_off_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( io_off_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( io_off_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( io_off_mem_rep_tag ),
       .mainOff_lock_req_ready( io_off_lock_req_ready ),
       .mainOff_lock_req_valid( mainComp_mainOff_lock_req_valid ),
       .mainOff_lock_req_bits_id(  ),
       .mainOff_lock_req_bits_op(  ),
       .mainOff_lock_req_tag( mainComp_mainOff_lock_req_tag ),
       .mainOff_lock_rep_ready( mainComp_mainOff_lock_rep_ready ),
       .mainOff_lock_rep_valid( io_off_lock_rep_valid ),
       .mainOff_lock_rep_bits_out(  ),
       .mainOff_lock_rep_tag( io_off_lock_rep_tag ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_7 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gRRDistributor_1(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_done,
    output[31:0] io_out_0_bits_pageId,
    output[63:0] io_out_0_bits_rankUpdate,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_done,
    output[31:0] io_out_1_bits_pageId,
    output[63:0] io_out_1_bits_rankUpdate,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output io_out_2_bits_done,
    output[31:0] io_out_2_bits_pageId,
    output[63:0] io_out_2_bits_rankUpdate,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output io_out_3_bits_done,
    output[31:0] io_out_3_bits_pageId,
    output[63:0] io_out_3_bits_rankUpdate,
    output[9:0] io_out_3_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    output[1:0] io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg[1:0] last_grant;
  wire T11;
  wire[1:0] T12;
  wire[1:0] choose;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;

  assign io_in_ready = T0;
  assign T0 = T73 || io_out_3_ready;
  assign io_out_1_valid = T1;
  assign T1 = T2 && io_in_valid;
  assign T2 = T55 || T3;
  assign T3 = ! T4;
  assign T4 = T52 || io_out_0_ready;
  assign io_out_0_valid = T5;
  assign T5 = T6 && io_in_valid;
  assign T6 = T50 || T7;
  assign T7 = ! T8;
  assign T8 = T48 || T9;
  assign T9 = io_out_3_ready && T10;
  assign T10 = 2'h3/* 3*/ > last_grant;
  assign T11 = io_in_valid && io_in_ready;
  assign T12 = T11 ? choose : last_grant;
  assign choose = T45 ? T44 : T13;
  assign T13 = T42 ? 2'h2/* 2*/ : T14;
  assign T14 = T40 ? 2'h3/* 3*/ : T15;
  assign T15 = io_out_0_ready ? T39 : T16;
  assign T16 = io_out_1_ready ? T38 : T17;
  assign T17 = io_out_2_ready ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign io_out_2_valid = T18;
  assign T18 = T19 && io_in_valid;
  assign T19 = T34 || T20;
  assign T20 = ! T21;
  assign T21 = T22 || io_out_1_ready;
  assign T22 = T23 || io_out_0_ready;
  assign T23 = T24 || T9;
  assign T24 = T27 || T25;
  assign T25 = io_out_2_ready && T26;
  assign T26 = 2'h2/* 2*/ > last_grant;
  assign T27 = T31 || T28;
  assign T28 = io_out_1_ready && T29;
  assign T29 = T30 > last_grant;
  assign T30 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T31 = io_out_0_ready && T32;
  assign T32 = T33 > last_grant;
  assign T33 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T34 = T36 && T35;
  assign T35 = 2'h2/* 2*/ > last_grant;
  assign T36 = ! T37;
  assign T37 = T31 || T28;
  assign io_out_2_bits_done = io_in_bits_done;
  assign T38 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T39 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T40 = io_out_3_ready && T41;
  assign T41 = 2'h3/* 3*/ > last_grant;
  assign T42 = io_out_2_ready && T43;
  assign T43 = 2'h2/* 2*/ > last_grant;
  assign T44 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T45 = io_out_1_ready && T46;
  assign T46 = T47 > last_grant;
  assign T47 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T48 = T49 || T25;
  assign T49 = T31 || T28;
  assign T50 = T51 > last_grant;
  assign T51 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign io_out_0_bits_done = io_in_bits_done;
  assign T52 = T53 || T9;
  assign T53 = T54 || T25;
  assign T54 = T31 || T28;
  assign T55 = T58 && T56;
  assign T56 = T57 > last_grant;
  assign T57 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T58 = ! T31;
  assign io_out_1_bits_done = io_in_bits_done;
  assign io_out_3_valid = T59;
  assign T59 = T60 && io_in_valid;
  assign T60 = T68 || T61;
  assign T61 = ! T62;
  assign T62 = T63 || io_out_2_ready;
  assign T63 = T64 || io_out_1_ready;
  assign T64 = T65 || io_out_0_ready;
  assign T65 = T66 || T9;
  assign T66 = T67 || T25;
  assign T67 = T31 || T28;
  assign T68 = T70 && T69;
  assign T69 = 2'h3/* 3*/ > last_grant;
  assign T70 = ! T71;
  assign T71 = T72 || T25;
  assign T72 = T31 || T28;
  assign io_out_3_bits_done = io_in_bits_done;
  assign io_out_2_bits_pageId = io_in_bits_pageId;
  assign io_out_1_bits_pageId = io_in_bits_pageId;
  assign io_out_0_bits_pageId = io_in_bits_pageId;
  assign io_out_3_bits_pageId = io_in_bits_pageId;
  assign T73 = T74 || io_out_2_ready;
  assign T74 = io_out_0_ready || io_out_1_ready;
  assign io_out_3_tag = io_in_tag;
  assign io_out_2_tag = io_in_tag;
  assign io_out_1_tag = io_in_tag;
  assign io_out_0_tag = io_in_tag;
  assign io_out_0_bits_rankUpdate = io_in_bits_rankUpdate;
  assign io_out_1_bits_rankUpdate = io_in_bits_rankUpdate;
  assign io_out_2_bits_rankUpdate = io_in_bits_rankUpdate;
  assign io_out_3_bits_rankUpdate = io_in_bits_rankUpdate;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T11) begin
      last_grant <= T12;
    end
  end
endmodule

module RRDistributorComponent_1(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_done,
    output[31:0] io_out_0_bits_pageId,
    output[63:0] io_out_0_bits_rankUpdate,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_done,
    output[31:0] io_out_1_bits_pageId,
    output[63:0] io_out_1_bits_rankUpdate,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output io_out_2_bits_done,
    output[31:0] io_out_2_bits_pageId,
    output[63:0] io_out_2_bits_rankUpdate,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output io_out_3_bits_done,
    output[31:0] io_out_3_bits_pageId,
    output[63:0] io_out_3_bits_rankUpdate,
    output[9:0] io_out_3_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    output[1:0] io_chosen);

  wire rrDist_io_in_ready;
  wire rrDist_io_out_1_valid;
  wire rrDist_io_out_0_valid;
  wire rrDist_io_out_2_valid;
  wire rrDist_io_out_2_bits_done;
  wire rrDist_io_out_0_bits_done;
  wire rrDist_io_out_1_bits_done;
  wire rrDist_io_out_3_valid;
  wire rrDist_io_out_3_bits_done;
  wire[31:0] rrDist_io_out_2_bits_pageId;
  wire[31:0] rrDist_io_out_1_bits_pageId;
  wire[31:0] rrDist_io_out_0_bits_pageId;
  wire[31:0] rrDist_io_out_3_bits_pageId;
  wire[9:0] rrDist_io_out_3_tag;
  wire[9:0] rrDist_io_out_2_tag;
  wire[9:0] rrDist_io_out_1_tag;
  wire[9:0] rrDist_io_out_0_tag;
  wire[63:0] rrDist_io_out_0_bits_rankUpdate;
  wire[63:0] rrDist_io_out_1_bits_rankUpdate;
  wire[63:0] rrDist_io_out_2_bits_rankUpdate;
  wire[63:0] rrDist_io_out_3_bits_rankUpdate;

  assign io_in_ready = rrDist_io_in_ready;
  assign io_out_1_valid = rrDist_io_out_1_valid;
  assign io_out_0_valid = rrDist_io_out_0_valid;
  assign io_out_2_valid = rrDist_io_out_2_valid;
  assign io_out_2_bits_done = rrDist_io_out_2_bits_done;
  assign io_out_0_bits_done = rrDist_io_out_0_bits_done;
  assign io_out_1_bits_done = rrDist_io_out_1_bits_done;
  assign io_out_3_valid = rrDist_io_out_3_valid;
  assign io_out_3_bits_done = rrDist_io_out_3_bits_done;
  assign io_out_2_bits_pageId = rrDist_io_out_2_bits_pageId;
  assign io_out_1_bits_pageId = rrDist_io_out_1_bits_pageId;
  assign io_out_0_bits_pageId = rrDist_io_out_0_bits_pageId;
  assign io_out_3_bits_pageId = rrDist_io_out_3_bits_pageId;
  assign io_out_3_tag = rrDist_io_out_3_tag;
  assign io_out_2_tag = rrDist_io_out_2_tag;
  assign io_out_1_tag = rrDist_io_out_1_tag;
  assign io_out_0_tag = rrDist_io_out_0_tag;
  assign io_out_0_bits_rankUpdate = rrDist_io_out_0_bits_rankUpdate;
  assign io_out_1_bits_rankUpdate = rrDist_io_out_1_bits_rankUpdate;
  assign io_out_2_bits_rankUpdate = rrDist_io_out_2_bits_rankUpdate;
  assign io_out_3_bits_rankUpdate = rrDist_io_out_3_bits_rankUpdate;
  gRRDistributor_1 rrDist(.clk(clk), .reset(reset),
       .io_out_0_ready( io_out_0_ready ),
       .io_out_0_valid( rrDist_io_out_0_valid ),
       .io_out_0_bits_done( rrDist_io_out_0_bits_done ),
       .io_out_0_bits_pageId( rrDist_io_out_0_bits_pageId ),
       .io_out_0_bits_rankUpdate( rrDist_io_out_0_bits_rankUpdate ),
       .io_out_0_tag( rrDist_io_out_0_tag ),
       .io_out_1_ready( io_out_1_ready ),
       .io_out_1_valid( rrDist_io_out_1_valid ),
       .io_out_1_bits_done( rrDist_io_out_1_bits_done ),
       .io_out_1_bits_pageId( rrDist_io_out_1_bits_pageId ),
       .io_out_1_bits_rankUpdate( rrDist_io_out_1_bits_rankUpdate ),
       .io_out_1_tag( rrDist_io_out_1_tag ),
       .io_out_2_ready( io_out_2_ready ),
       .io_out_2_valid( rrDist_io_out_2_valid ),
       .io_out_2_bits_done( rrDist_io_out_2_bits_done ),
       .io_out_2_bits_pageId( rrDist_io_out_2_bits_pageId ),
       .io_out_2_bits_rankUpdate( rrDist_io_out_2_bits_rankUpdate ),
       .io_out_2_tag( rrDist_io_out_2_tag ),
       .io_out_3_ready( io_out_3_ready ),
       .io_out_3_valid( rrDist_io_out_3_valid ),
       .io_out_3_bits_done( rrDist_io_out_3_bits_done ),
       .io_out_3_bits_pageId( rrDist_io_out_3_bits_pageId ),
       .io_out_3_bits_rankUpdate( rrDist_io_out_3_bits_rankUpdate ),
       .io_out_3_tag( rrDist_io_out_3_tag ),
       .io_in_ready( rrDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
endmodule

module gRRArbiter_1(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_out,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_out,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_out,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_out,
    input [9:0] io_in_3_tag,
    output[1:0] io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire[1:0] choose;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[9:0] T75;
  wire[4:0] T76;
  wire[4:0] T77;
  wire[4:0] T78;
  wire T79;
  wire[3:0] T80;
  wire[6:0] T81;
  wire[4:0] tvec_3;
  wire[4:0] T82;
  wire[4:0] T83;
  wire[4:0] T84;
  wire[4:0] T85;
  wire T86;
  wire[4:0] tvec_2;
  wire[4:0] T87;
  wire[4:0] T88;
  wire[4:0] T89;
  wire[4:0] T90;
  wire T91;
  wire[4:0] tvec_1;
  wire[4:0] T92;
  wire[4:0] T93;
  wire[4:0] T94;
  wire T95;
  wire[4:0] tvec_0;
  wire[4:0] T96;

  assign io_in_2_ready = T0;
  assign T0 = T1 && io_out_ready;
  assign T1 = T38 || T2;
  assign T2 = ! T3;
  assign T3 = T4 || io_in_1_valid;
  assign T4 = T5 || io_in_0_valid;
  assign T5 = T28 || T6;
  assign T6 = io_in_3_valid && T7;
  assign T7 = 2'h3/* 3*/ > last_grant;
  assign T8 = io_out_valid && io_out_ready;
  assign io_out_valid = T9;
  assign T9 = T10 || io_in_3_valid;
  assign T10 = T11 || io_in_2_valid;
  assign T11 = io_in_0_valid || io_in_1_valid;
  assign T12 = T8 ? choose : last_grant;
  assign choose = T25 ? T24 : T13;
  assign T13 = T22 ? 2'h2/* 2*/ : T14;
  assign T14 = T20 ? 2'h3/* 3*/ : T15;
  assign T15 = io_in_0_valid ? T19 : T16;
  assign T16 = io_in_1_valid ? T18 : T17;
  assign T17 = io_in_2_valid ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T18 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T19 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T20 = io_in_3_valid && T21;
  assign T21 = 2'h3/* 3*/ > last_grant;
  assign T22 = io_in_2_valid && T23;
  assign T23 = 2'h2/* 2*/ > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T25 = io_in_1_valid && T26;
  assign T26 = T27 > last_grant;
  assign T27 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T28 = T31 || T29;
  assign T29 = io_in_2_valid && T30;
  assign T30 = 2'h2/* 2*/ > last_grant;
  assign T31 = T35 || T32;
  assign T32 = io_in_1_valid && T33;
  assign T33 = T34 > last_grant;
  assign T34 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T35 = io_in_0_valid && T36;
  assign T36 = T37 > last_grant;
  assign T37 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T38 = T40 && T39;
  assign T39 = 2'h2/* 2*/ > last_grant;
  assign T40 = ! T41;
  assign T41 = T35 || T32;
  assign io_in_0_ready = T42;
  assign T42 = T43 && io_out_ready;
  assign T43 = T48 || T44;
  assign T44 = ! T45;
  assign T45 = T46 || T6;
  assign T46 = T47 || T29;
  assign T47 = T35 || T32;
  assign T48 = T49 > last_grant;
  assign T49 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign io_in_1_ready = T50;
  assign T50 = T51 && io_out_ready;
  assign T51 = T57 || T52;
  assign T52 = ! T53;
  assign T53 = T54 || io_in_0_valid;
  assign T54 = T55 || T6;
  assign T55 = T56 || T29;
  assign T56 = T35 || T32;
  assign T57 = T60 && T58;
  assign T58 = T59 > last_grant;
  assign T59 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T60 = ! T35;
  assign io_in_3_ready = T61;
  assign T61 = T62 && io_out_ready;
  assign T62 = T70 || T63;
  assign T63 = ! T64;
  assign T64 = T65 || io_in_2_valid;
  assign T65 = T66 || io_in_1_valid;
  assign T66 = T67 || io_in_0_valid;
  assign T67 = T68 || T6;
  assign T68 = T69 || T29;
  assign T69 = T35 || T32;
  assign T70 = T72 && T71;
  assign T71 = 2'h3/* 3*/ > last_grant;
  assign T72 = ! T73;
  assign T73 = T74 || T29;
  assign T74 = T35 || T32;
  assign io_out_tag = T75;
  assign T75 = {5'h0/* 0*/, T76};
  assign T76 = T83 | T77;
  assign T77 = tvec_3 & T78;
  assign T78 = {3'h5/* 5*/{T79}};
  assign T79 = T80[2'h3/* 3*/];
  assign T80 = T81[2'h3/* 3*/:1'h0/* 0*/];
  assign T81 = 4'h1/* 1*/ << choose;
  assign tvec_3 = T82;
  assign T82 = io_in_3_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T83 = T88 | T84;
  assign T84 = tvec_2 & T85;
  assign T85 = {3'h5/* 5*/{T86}};
  assign T86 = T80[2'h2/* 2*/];
  assign tvec_2 = T87;
  assign T87 = io_in_2_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T88 = T93 | T89;
  assign T89 = tvec_1 & T90;
  assign T90 = {3'h5/* 5*/{T91}};
  assign T91 = T80[1'h1/* 1*/];
  assign tvec_1 = T92;
  assign T92 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T93 = tvec_0 & T94;
  assign T94 = {3'h5/* 5*/{T95}};
  assign T95 = T80[1'h0/* 0*/];
  assign tvec_0 = T96;
  assign T96 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T12;
    end
  end
endmodule

module RRAggregatorComponent_1(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_out,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_out,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_out,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_out,
    input [9:0] io_in_3_tag,
    output[1:0] io_chosen);

  wire rrArb_io_in_2_ready;
  wire rrArb_io_in_0_ready;
  wire rrArb_io_in_1_ready;
  wire rrArb_io_in_3_ready;
  wire[9:0] rrArb_io_out_tag;
  wire rrArb_io_out_valid;

  assign io_in_2_ready = rrArb_io_in_2_ready;
  assign io_in_0_ready = rrArb_io_in_0_ready;
  assign io_in_1_ready = rrArb_io_in_1_ready;
  assign io_in_3_ready = rrArb_io_in_3_ready;
  assign io_out_tag = rrArb_io_out_tag;
  assign io_out_valid = rrArb_io_out_valid;
  gRRArbiter_1 rrArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( rrArb_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( rrArb_io_out_tag ),
       .io_in_0_ready( rrArb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_valid ),
       .io_in_0_bits_out(  ),
       .io_in_0_tag( io_in_0_tag ),
       .io_in_1_ready( rrArb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_valid ),
       .io_in_1_bits_out(  ),
       .io_in_1_tag( io_in_1_tag ),
       .io_in_2_ready( rrArb_io_in_2_ready ),
       .io_in_2_valid( io_in_2_valid ),
       .io_in_2_bits_out(  ),
       .io_in_2_tag( io_in_2_tag ),
       .io_in_3_ready( rrArb_io_in_3_ready ),
       .io_in_3_valid( io_in_3_valid ),
       .io_in_3_bits_out(  ),
       .io_in_3_tag( io_in_3_tag ),
       .io_chosen(  ));
endmodule

module gTaggedRRArbiter_1(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_addr,
    output io_out_bits_rw,
    output io_out_bits_cached,
    output[127:0] io_out_bits_data,
    output[3:0] io_out_bits_size,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_addr,
    input  io_in_0_bits_rw,
    input  io_in_0_bits_cached,
    input [127:0] io_in_0_bits_data,
    input [3:0] io_in_0_bits_size,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_addr,
    input  io_in_1_bits_rw,
    input  io_in_1_bits_cached,
    input [127:0] io_in_1_bits_data,
    input [3:0] io_in_1_bits_size,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [31:0] io_in_2_bits_addr,
    input  io_in_2_bits_rw,
    input  io_in_2_bits_cached,
    input [127:0] io_in_2_bits_data,
    input [3:0] io_in_2_bits_size,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [31:0] io_in_3_bits_addr,
    input  io_in_3_bits_rw,
    input  io_in_3_bits_cached,
    input [127:0] io_in_3_bits_data,
    input [3:0] io_in_3_bits_size,
    input [9:0] io_in_3_tag,
    output[1:0] io_chosen);

  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire T3;
  wire[3:0] T4;
  wire[6:0] T5;
  wire[1:0] choose;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg[1:0] last_grant;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[1:0] T66;
  wire[3:0] dvec_3_size;
  wire[31:0] T67;
  wire[31:0] T68;
  wire[31:0] T69;
  wire[31:0] dvec_3_addr;
  wire[31:0] T70;
  wire[31:0] T71;
  wire[31:0] T72;
  wire T73;
  wire[31:0] dvec_2_addr;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[31:0] T76;
  wire T77;
  wire[31:0] dvec_1_addr;
  wire[31:0] T78;
  wire[31:0] T79;
  wire T80;
  wire[31:0] dvec_0_addr;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire[3:0] dvec_2_size;
  wire[3:0] T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire[3:0] dvec_1_size;
  wire[3:0] T87;
  wire[3:0] T88;
  wire[3:0] dvec_0_size;
  wire[127:0] T89;
  wire[127:0] T90;
  wire[127:0] T91;
  wire[127:0] dvec_3_data;
  wire[127:0] T92;
  wire[127:0] T93;
  wire[127:0] T94;
  wire[127:0] dvec_2_data;
  wire[127:0] T95;
  wire[127:0] T96;
  wire[127:0] T97;
  wire[127:0] dvec_1_data;
  wire[127:0] T98;
  wire[127:0] T99;
  wire[127:0] dvec_0_data;
  wire T100;
  wire T101;
  wire dvec_3_cached;
  wire T102;
  wire T103;
  wire dvec_2_cached;
  wire T104;
  wire T105;
  wire dvec_1_cached;
  wire T106;
  wire dvec_0_cached;
  wire T107;
  wire T108;
  wire dvec_3_rw;
  wire T109;
  wire T110;
  wire dvec_2_rw;
  wire T111;
  wire T112;
  wire dvec_1_rw;
  wire T113;
  wire dvec_0_rw;
  wire[9:0] T114;
  wire[6:0] T115;
  wire[6:0] T116;
  wire[6:0] T117;
  wire[4:0] T118;
  wire[4:0] T119;
  wire[4:0] T120;
  wire[4:0] tvec_3;
  wire[4:0] T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire[4:0] T124;
  wire[4:0] tvec_2;
  wire[4:0] T125;
  wire[4:0] T126;
  wire[4:0] T127;
  wire[4:0] T128;
  wire[4:0] tvec_1;
  wire[4:0] T129;
  wire[4:0] T130;
  wire[4:0] T131;
  wire[4:0] tvec_0;
  wire[4:0] T132;
  wire[6:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;

  assign io_out_bits_size = T0;
  assign T0 = T81 | T1;
  assign T1 = dvec_3_size & T2;
  assign T2 = {3'h4/* 4*/{T3}};
  assign T3 = T4[2'h3/* 3*/];
  assign T4 = T5[2'h3/* 3*/:1'h0/* 0*/];
  assign T5 = 4'h1/* 1*/ << choose;
  assign choose = T64 ? T63 : T6;
  assign T6 = T61 ? 2'h2/* 2*/ : T7;
  assign T7 = T59 ? 2'h3/* 3*/ : T8;
  assign T8 = io_in_0_valid ? T58 : T9;
  assign T9 = io_in_1_valid ? T11 : T10;
  assign T10 = io_in_2_valid ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign io_in_0_ready = T12;
  assign T12 = T13 && io_out_ready;
  assign T13 = T33 || T14;
  assign T14 = ! T15;
  assign T15 = T23 || T16;
  assign T16 = io_in_3_valid && T17;
  assign T17 = 2'h3/* 3*/ > last_grant;
  assign T18 = io_out_valid && io_out_ready;
  assign io_out_valid = T19;
  assign T19 = T20 || io_in_3_valid;
  assign T20 = T21 || io_in_2_valid;
  assign T21 = io_in_0_valid || io_in_1_valid;
  assign T22 = T18 ? choose : last_grant;
  assign T23 = T26 || T24;
  assign T24 = io_in_2_valid && T25;
  assign T25 = 2'h2/* 2*/ > last_grant;
  assign T26 = T30 || T27;
  assign T27 = io_in_1_valid && T28;
  assign T28 = T29 > last_grant;
  assign T29 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T30 = io_in_0_valid && T31;
  assign T31 = T32 > last_grant;
  assign T32 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T33 = T34 > last_grant;
  assign T34 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign io_in_2_ready = T35;
  assign T35 = T36 && io_out_ready;
  assign T36 = T43 || T37;
  assign T37 = ! T38;
  assign T38 = T39 || io_in_1_valid;
  assign T39 = T40 || io_in_0_valid;
  assign T40 = T41 || T16;
  assign T41 = T42 || T24;
  assign T42 = T30 || T27;
  assign T43 = T45 && T44;
  assign T44 = 2'h2/* 2*/ > last_grant;
  assign T45 = ! T46;
  assign T46 = T30 || T27;
  assign io_in_1_ready = T47;
  assign T47 = T48 && io_out_ready;
  assign T48 = T54 || T49;
  assign T49 = ! T50;
  assign T50 = T51 || io_in_0_valid;
  assign T51 = T52 || T16;
  assign T52 = T53 || T24;
  assign T53 = T30 || T27;
  assign T54 = T57 && T55;
  assign T55 = T56 > last_grant;
  assign T56 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T57 = ! T30;
  assign T58 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T59 = io_in_3_valid && T60;
  assign T60 = 2'h3/* 3*/ > last_grant;
  assign T61 = io_in_2_valid && T62;
  assign T62 = 2'h2/* 2*/ > last_grant;
  assign T63 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T64 = io_in_1_valid && T65;
  assign T65 = T66 > last_grant;
  assign T66 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign dvec_3_size = io_in_3_bits_size;
  assign io_out_bits_addr = T67;
  assign T67 = T70 | T68;
  assign T68 = dvec_3_addr & T69;
  assign T69 = {6'h20/* 32*/{T3}};
  assign dvec_3_addr = io_in_3_bits_addr;
  assign T70 = T74 | T71;
  assign T71 = dvec_2_addr & T72;
  assign T72 = {6'h20/* 32*/{T73}};
  assign T73 = T4[2'h2/* 2*/];
  assign dvec_2_addr = io_in_2_bits_addr;
  assign T74 = T78 | T75;
  assign T75 = dvec_1_addr & T76;
  assign T76 = {6'h20/* 32*/{T77}};
  assign T77 = T4[1'h1/* 1*/];
  assign dvec_1_addr = io_in_1_bits_addr;
  assign T78 = dvec_0_addr & T79;
  assign T79 = {6'h20/* 32*/{T80}};
  assign T80 = T4[1'h0/* 0*/];
  assign dvec_0_addr = io_in_0_bits_addr;
  assign T81 = T84 | T82;
  assign T82 = dvec_2_size & T83;
  assign T83 = {3'h4/* 4*/{T73}};
  assign dvec_2_size = io_in_2_bits_size;
  assign T84 = T87 | T85;
  assign T85 = dvec_1_size & T86;
  assign T86 = {3'h4/* 4*/{T77}};
  assign dvec_1_size = io_in_1_bits_size;
  assign T87 = dvec_0_size & T88;
  assign T88 = {3'h4/* 4*/{T80}};
  assign dvec_0_size = io_in_0_bits_size;
  assign io_out_bits_data = T89;
  assign T89 = T92 | T90;
  assign T90 = dvec_3_data & T91;
  assign T91 = {8'h80/* 128*/{T3}};
  assign dvec_3_data = io_in_3_bits_data;
  assign T92 = T95 | T93;
  assign T93 = dvec_2_data & T94;
  assign T94 = {8'h80/* 128*/{T73}};
  assign dvec_2_data = io_in_2_bits_data;
  assign T95 = T98 | T96;
  assign T96 = dvec_1_data & T97;
  assign T97 = {8'h80/* 128*/{T77}};
  assign dvec_1_data = io_in_1_bits_data;
  assign T98 = dvec_0_data & T99;
  assign T99 = {8'h80/* 128*/{T80}};
  assign dvec_0_data = io_in_0_bits_data;
  assign io_out_bits_cached = T100;
  assign T100 = T102 | T101;
  assign T101 = dvec_3_cached & T3;
  assign dvec_3_cached = io_in_3_bits_cached;
  assign T102 = T104 | T103;
  assign T103 = dvec_2_cached & T73;
  assign dvec_2_cached = io_in_2_bits_cached;
  assign T104 = T106 | T105;
  assign T105 = dvec_1_cached & T77;
  assign dvec_1_cached = io_in_1_bits_cached;
  assign T106 = dvec_0_cached & T80;
  assign dvec_0_cached = io_in_0_bits_cached;
  assign io_out_bits_rw = T107;
  assign T107 = T109 | T108;
  assign T108 = dvec_3_rw & T3;
  assign dvec_3_rw = io_in_3_bits_rw;
  assign T109 = T111 | T110;
  assign T110 = dvec_2_rw & T73;
  assign dvec_2_rw = io_in_2_bits_rw;
  assign T111 = T113 | T112;
  assign T112 = dvec_1_rw & T77;
  assign dvec_1_rw = io_in_1_bits_rw;
  assign T113 = dvec_0_rw & T80;
  assign dvec_0_rw = io_in_0_bits_rw;
  assign io_out_tag = T114;
  assign T114 = {3'h0/* 0*/, T115};
  assign T115 = T133 | T116;
  assign T116 = T117 & 7'h1f/* 31*/;
  assign T117 = {2'h0/* 0*/, T118};
  assign T118 = T122 | T119;
  assign T119 = tvec_3 & T120;
  assign T120 = {3'h5/* 5*/{T3}};
  assign tvec_3 = T121;
  assign T121 = io_in_3_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T122 = T126 | T123;
  assign T123 = tvec_2 & T124;
  assign T124 = {3'h5/* 5*/{T73}};
  assign tvec_2 = T125;
  assign T125 = io_in_2_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T126 = T130 | T127;
  assign T127 = tvec_1 & T128;
  assign T128 = {3'h5/* 5*/{T77}};
  assign tvec_1 = T129;
  assign T129 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T130 = tvec_0 & T131;
  assign T131 = {3'h5/* 5*/{T80}};
  assign tvec_0 = T132;
  assign T132 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T133 = choose << 3'h5/* 5*/;
  assign io_in_3_ready = T134;
  assign T134 = T135 && io_out_ready;
  assign T135 = T143 || T136;
  assign T136 = ! T137;
  assign T137 = T138 || io_in_2_valid;
  assign T138 = T139 || io_in_1_valid;
  assign T139 = T140 || io_in_0_valid;
  assign T140 = T141 || T16;
  assign T141 = T142 || T24;
  assign T142 = T30 || T27;
  assign T143 = T145 && T144;
  assign T144 = 2'h3/* 3*/ > last_grant;
  assign T145 = ! T146;
  assign T146 = T147 || T24;
  assign T147 = T30 || T27;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T18) begin
      last_grant <= T22;
    end
  end
endmodule

module gTaggedRRArbiter_2(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_id,
    output io_out_bits_op,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_id,
    input  io_in_0_bits_op,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_id,
    input  io_in_1_bits_op,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [31:0] io_in_2_bits_id,
    input  io_in_2_bits_op,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [31:0] io_in_3_bits_id,
    input  io_in_3_bits_op,
    input [9:0] io_in_3_tag,
    output[1:0] io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire[1:0] T9;
  wire[1:0] choose;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[1:0] T31;
  wire T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire[9:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire[4:0] T65;
  wire[4:0] T66;
  wire[4:0] T67;
  wire T68;
  wire[3:0] T69;
  wire[6:0] T70;
  wire[4:0] tvec_3;
  wire[4:0] T71;
  wire[4:0] T72;
  wire[4:0] T73;
  wire[4:0] T74;
  wire T75;
  wire[4:0] tvec_2;
  wire[4:0] T76;
  wire[4:0] T77;
  wire[4:0] T78;
  wire[4:0] T79;
  wire T80;
  wire[4:0] tvec_1;
  wire[4:0] T81;
  wire[4:0] T82;
  wire[4:0] T83;
  wire T84;
  wire[4:0] tvec_0;
  wire[4:0] T85;
  wire[6:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;

  assign io_out_valid = T0;
  assign T0 = T1 || io_in_3_valid;
  assign T1 = T60 || io_in_2_valid;
  assign io_in_0_ready = T2;
  assign T2 = T3 && io_out_ready;
  assign T3 = T35 || T4;
  assign T4 = ! T5;
  assign T5 = T25 || T6;
  assign T6 = io_in_3_valid && T7;
  assign T7 = 2'h3/* 3*/ > last_grant;
  assign T8 = io_out_valid && io_out_ready;
  assign T9 = T8 ? choose : last_grant;
  assign choose = T22 ? T21 : T10;
  assign T10 = T19 ? 2'h2/* 2*/ : T11;
  assign T11 = T17 ? 2'h3/* 3*/ : T12;
  assign T12 = io_in_0_valid ? T16 : T13;
  assign T13 = io_in_1_valid ? T15 : T14;
  assign T14 = io_in_2_valid ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T15 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T16 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T17 = io_in_3_valid && T18;
  assign T18 = 2'h3/* 3*/ > last_grant;
  assign T19 = io_in_2_valid && T20;
  assign T20 = 2'h2/* 2*/ > last_grant;
  assign T21 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T22 = io_in_1_valid && T23;
  assign T23 = T24 > last_grant;
  assign T24 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T25 = T28 || T26;
  assign T26 = io_in_2_valid && T27;
  assign T27 = 2'h2/* 2*/ > last_grant;
  assign T28 = T32 || T29;
  assign T29 = io_in_1_valid && T30;
  assign T30 = T31 > last_grant;
  assign T31 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T32 = io_in_0_valid && T33;
  assign T33 = T34 > last_grant;
  assign T34 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T35 = T36 > last_grant;
  assign T36 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign io_in_2_ready = T37;
  assign T37 = T38 && io_out_ready;
  assign T38 = T45 || T39;
  assign T39 = ! T40;
  assign T40 = T41 || io_in_1_valid;
  assign T41 = T42 || io_in_0_valid;
  assign T42 = T43 || T6;
  assign T43 = T44 || T26;
  assign T44 = T32 || T29;
  assign T45 = T47 && T46;
  assign T46 = 2'h2/* 2*/ > last_grant;
  assign T47 = ! T48;
  assign T48 = T32 || T29;
  assign io_in_1_ready = T49;
  assign T49 = T50 && io_out_ready;
  assign T50 = T56 || T51;
  assign T51 = ! T52;
  assign T52 = T53 || io_in_0_valid;
  assign T53 = T54 || T6;
  assign T54 = T55 || T26;
  assign T55 = T32 || T29;
  assign T56 = T59 && T57;
  assign T57 = T58 > last_grant;
  assign T58 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T59 = ! T32;
  assign T60 = io_in_0_valid || io_in_1_valid;
  assign io_out_tag = T61;
  assign T61 = {3'h0/* 0*/, T62};
  assign T62 = T86 | T63;
  assign T63 = T64 & 7'h1f/* 31*/;
  assign T64 = {2'h0/* 0*/, T65};
  assign T65 = T72 | T66;
  assign T66 = tvec_3 & T67;
  assign T67 = {3'h5/* 5*/{T68}};
  assign T68 = T69[2'h3/* 3*/];
  assign T69 = T70[2'h3/* 3*/:1'h0/* 0*/];
  assign T70 = 4'h1/* 1*/ << choose;
  assign tvec_3 = T71;
  assign T71 = io_in_3_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T72 = T77 | T73;
  assign T73 = tvec_2 & T74;
  assign T74 = {3'h5/* 5*/{T75}};
  assign T75 = T69[2'h2/* 2*/];
  assign tvec_2 = T76;
  assign T76 = io_in_2_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T77 = T82 | T78;
  assign T78 = tvec_1 & T79;
  assign T79 = {3'h5/* 5*/{T80}};
  assign T80 = T69[1'h1/* 1*/];
  assign tvec_1 = T81;
  assign T81 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T82 = tvec_0 & T83;
  assign T83 = {3'h5/* 5*/{T84}};
  assign T84 = T69[1'h0/* 0*/];
  assign tvec_0 = T85;
  assign T85 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T86 = choose << 3'h5/* 5*/;
  assign io_in_3_ready = T87;
  assign T87 = T88 && io_out_ready;
  assign T88 = T96 || T89;
  assign T89 = ! T90;
  assign T90 = T91 || io_in_2_valid;
  assign T91 = T92 || io_in_1_valid;
  assign T92 = T93 || io_in_0_valid;
  assign T93 = T94 || T6;
  assign T94 = T95 || T26;
  assign T95 = T32 || T29;
  assign T96 = T98 && T97;
  assign T97 = 2'h3/* 3*/ > last_grant;
  assign T98 = ! T99;
  assign T99 = T100 || T26;
  assign T100 = T32 || T29;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T9;
    end
  end
endmodule

module gTaggedDistributor_1(
    input  io_out_0_ready,
    output io_out_0_valid,
    output[127:0] io_out_0_bits_data,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[127:0] io_out_1_bits_data,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[127:0] io_out_2_bits_data,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output[127:0] io_out_3_bits_data,
    output[9:0] io_out_3_tag,
    output io_in_ready,
    input  io_in_valid,
    input [127:0] io_in_bits_data,
    input [9:0] io_in_tag,
    output[1:0] io_chosen);

  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T2;
  wire[9:0] T3;
  wire T4;
  wire T5;
  wire[9:0] T6;
  wire[9:0] T7;
  wire[9:0] T8;
  wire[9:0] T9;
  wire[9:0] T10;
  wire[9:0] T11;
  wire T12;
  wire T13;
  wire[9:0] T14;
  wire[9:0] T15;
  wire[9:0] T16;
  wire[9:0] T17;
  wire[9:0] T18;
  wire[9:0] T19;
  wire T20;
  wire T21;
  wire[9:0] T22;
  wire[9:0] T23;
  wire[9:0] T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire[9:0] T28;
  wire[9:0] T29;
  wire[9:0] T30;
  wire[9:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire[1026:0] T37;
  wire[9:0] T38;
  wire[9:0] T39;
  wire[9:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;

  assign io_out_2_tag = T0;
  assign T0 = io_in_tag & T1;
  assign T1 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_1_tag = T2;
  assign T2 = io_in_tag & T3;
  assign T3 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_1_valid = T4;
  assign T4 = io_in_valid && T5;
  assign T5 = T9 == T6;
  assign T6 = T8 & T7;
  assign T7 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T8 = io_in_tag >> 3'h5/* 5*/;
  assign T9 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign io_out_0_tag = T10;
  assign T10 = io_in_tag & T11;
  assign T11 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_0_valid = T12;
  assign T12 = io_in_valid && T13;
  assign T13 = T17 == T14;
  assign T14 = T16 & T15;
  assign T15 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T16 = io_in_tag >> 3'h5/* 5*/;
  assign T17 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign io_out_3_tag = T18;
  assign T18 = io_in_tag & T19;
  assign T19 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_3_valid = T20;
  assign T20 = io_in_valid && T21;
  assign T21 = T25 == T22;
  assign T22 = T24 & T23;
  assign T23 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T24 = io_in_tag >> 3'h5/* 5*/;
  assign T25 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign io_out_3_bits_data = io_in_bits_data;
  assign io_out_2_valid = T26;
  assign T26 = io_in_valid && T27;
  assign T27 = T31 == T28;
  assign T28 = T30 & T29;
  assign T29 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T30 = io_in_tag >> 3'h5/* 5*/;
  assign T31 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign io_out_2_bits_data = io_in_bits_data;
  assign io_out_1_bits_data = io_in_bits_data;
  assign io_out_0_bits_data = io_in_bits_data;
  assign io_in_ready = T32;
  assign T32 = io_in_valid && T33;
  assign T33 = T41 | T34;
  assign T34 = io_out_3_ready & T35;
  assign T35 = T36[2'h3/* 3*/];
  assign T36 = T37[2'h3/* 3*/:1'h0/* 0*/];
  assign T37 = 4'h1/* 1*/ << T38;
  assign T38 = T40 & T39;
  assign T39 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T40 = io_in_tag >> 3'h5/* 5*/;
  assign T41 = T44 | T42;
  assign T42 = io_out_2_ready & T43;
  assign T43 = T36[2'h2/* 2*/];
  assign T44 = T47 | T45;
  assign T45 = io_out_1_ready & T46;
  assign T46 = T36[1'h1/* 1*/];
  assign T47 = io_out_0_ready & T48;
  assign T48 = T36[1'h0/* 0*/];
endmodule

module gTaggedDistributor_2(
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_out,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_out,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output io_out_2_bits_out,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output io_out_3_bits_out,
    output[9:0] io_out_3_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_out,
    input [9:0] io_in_tag,
    output[1:0] io_chosen);

  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T2;
  wire[9:0] T3;
  wire T4;
  wire T5;
  wire[9:0] T6;
  wire[9:0] T7;
  wire[9:0] T8;
  wire[9:0] T9;
  wire[9:0] T10;
  wire[9:0] T11;
  wire T12;
  wire T13;
  wire[9:0] T14;
  wire[9:0] T15;
  wire[9:0] T16;
  wire[9:0] T17;
  wire[9:0] T18;
  wire[9:0] T19;
  wire T20;
  wire T21;
  wire[9:0] T22;
  wire[9:0] T23;
  wire[9:0] T24;
  wire[9:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[3:0] T30;
  wire[1026:0] T31;
  wire[9:0] T32;
  wire[9:0] T33;
  wire[9:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[9:0] T45;
  wire[9:0] T46;
  wire[9:0] T47;
  wire[9:0] T48;

  assign io_out_3_tag = T0;
  assign T0 = io_in_tag & T1;
  assign T1 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_2_tag = T2;
  assign T2 = io_in_tag & T3;
  assign T3 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_2_valid = T4;
  assign T4 = io_in_valid && T5;
  assign T5 = T9 == T6;
  assign T6 = T8 & T7;
  assign T7 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T8 = io_in_tag >> 3'h5/* 5*/;
  assign T9 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign io_out_1_tag = T10;
  assign T10 = io_in_tag & T11;
  assign T11 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_1_valid = T12;
  assign T12 = io_in_valid && T13;
  assign T13 = T17 == T14;
  assign T14 = T16 & T15;
  assign T15 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T16 = io_in_tag >> 3'h5/* 5*/;
  assign T17 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign io_out_0_tag = T18;
  assign T18 = io_in_tag & T19;
  assign T19 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign io_out_0_valid = T20;
  assign T20 = io_in_valid && T21;
  assign T21 = T25 == T22;
  assign T22 = T24 & T23;
  assign T23 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T24 = io_in_tag >> 3'h5/* 5*/;
  assign T25 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign io_in_ready = T26;
  assign T26 = io_in_valid && T27;
  assign T27 = T35 | T28;
  assign T28 = io_out_3_ready & T29;
  assign T29 = T30[2'h3/* 3*/];
  assign T30 = T31[2'h3/* 3*/:1'h0/* 0*/];
  assign T31 = 4'h1/* 1*/ << T32;
  assign T32 = T34 & T33;
  assign T33 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T34 = io_in_tag >> 3'h5/* 5*/;
  assign T35 = T38 | T36;
  assign T36 = io_out_2_ready & T37;
  assign T37 = T30[2'h2/* 2*/];
  assign T38 = T41 | T39;
  assign T39 = io_out_1_ready & T40;
  assign T40 = T30[1'h1/* 1*/];
  assign T41 = io_out_0_ready & T42;
  assign T42 = T30[1'h0/* 0*/];
  assign io_out_3_valid = T43;
  assign T43 = io_in_valid && T44;
  assign T44 = T48 == T45;
  assign T45 = T47 & T46;
  assign T46 = {3'h0/* 0*/, 7'h1f/* 31*/};
  assign T47 = io_in_tag >> 3'h5/* 5*/;
  assign T48 = {5'h0/* 0*/, 5'h3/* 3*/};
endmodule

module gReplicatedComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag,
    input  mainOff_lock_req_ready,
    output mainOff_lock_req_valid,
    output[31:0] mainOff_lock_req_bits_id,
    output mainOff_lock_req_bits_op,
    output[9:0] mainOff_lock_req_tag,
    output mainOff_lock_rep_ready,
    input  mainOff_lock_rep_valid,
    input  mainOff_lock_rep_bits_out,
    input [9:0] mainOff_lock_rep_tag);

  wire inputDist_io_in_ready;
  wire gOffloadedComponent_3_io_in_ready;
  wire[9:0] gTaggedDistributor_1_io_out_3_tag;
  wire gTaggedRRArbiter_1_io_out_valid;
  wire gOffloadedComponent_3_io_off_lock_req_valid;
  wire gOffloadedComponent_2_io_off_lock_req_valid;
  wire[9:0] gTaggedDistributor_1_io_out_2_tag;
  wire gTaggedDistributor_1_io_out_2_valid;
  wire[9:0] gTaggedDistributor_io_out_2_tag;
  wire[3:0] gTaggedRRArbiter_io_out_bits_size;
  wire gOffloadedComponent_2_io_off_mem_req_valid;
  wire gOffloadedComponent_1_io_off_mem_req_valid;
  wire[9:0] gTaggedDistributor_1_io_out_1_tag;
  wire gTaggedDistributor_1_io_out_1_valid;
  wire[9:0] gTaggedDistributor_io_out_1_tag;
  wire gTaggedDistributor_io_out_1_valid;
  wire inputDist_io_out_1_valid;
  wire gOffloadedComponent_io_in_ready;
  wire[9:0] gTaggedDistributor_1_io_out_0_tag;
  wire gTaggedDistributor_1_io_out_0_valid;
  wire gTaggedRRArbiter_1_io_in_0_ready;
  wire gTaggedDistributor_1_io_in_ready;
  wire gOffloadedComponent_3_io_off_lock_rep_ready;
  wire gOffloadedComponent_2_io_off_lock_rep_ready;
  wire gOffloadedComponent_1_io_off_lock_rep_ready;
  wire gOffloadedComponent_io_off_lock_rep_ready;
  wire gOffloadedComponent_1_io_off_lock_req_valid;
  wire gOffloadedComponent_io_off_lock_req_valid;
  wire[9:0] gTaggedDistributor_io_out_0_tag;
  wire gTaggedDistributor_io_out_0_valid;
  wire gTaggedRRArbiter_io_in_0_ready;
  wire gOffloadedComponent_3_io_off_mem_req_valid;
  wire[9:0] gTaggedDistributor_io_out_3_tag;
  wire gTaggedDistributor_io_out_3_valid;
  wire gOffloadedComponent_io_off_mem_req_valid;
  wire inputDist_io_out_0_valid;
  wire gOffloadedComponent_2_io_in_ready;
  wire inputDist_io_out_2_valid;
  wire gOffloadedComponent_1_io_in_ready;
  wire inputDist_io_out_2_bits_done;
  wire outputArb_io_in_2_ready;
  wire gOffloadedComponent_1_io_out_valid;
  wire gOffloadedComponent_io_out_valid;
  wire gOffloadedComponent_3_io_out_valid;
  wire gOffloadedComponent_2_io_out_valid;
  wire gTaggedRRArbiter_1_io_in_2_ready;
  wire gTaggedRRArbiter_io_in_2_ready;
  wire inputDist_io_out_0_bits_done;
  wire outputArb_io_in_0_ready;
  wire inputDist_io_out_1_bits_done;
  wire outputArb_io_in_1_ready;
  wire gTaggedRRArbiter_1_io_in_1_ready;
  wire gTaggedRRArbiter_io_in_1_ready;
  wire[3:0] gOffloadedComponent_3_io_off_mem_req_bits_size;
  wire inputDist_io_out_3_valid;
  wire inputDist_io_out_3_bits_done;
  wire outputArb_io_in_3_ready;
  wire[127:0] gTaggedDistributor_io_out_3_bits_data;
  wire[31:0] gTaggedRRArbiter_io_out_bits_addr;
  wire[31:0] gOffloadedComponent_3_io_off_mem_req_bits_addr;
  wire[31:0] gOffloadedComponent_2_io_off_mem_req_bits_addr;
  wire gTaggedDistributor_io_out_2_valid;
  wire[127:0] gTaggedDistributor_io_out_2_bits_data;
  wire[31:0] inputDist_io_out_2_bits_pageId;
  wire[31:0] gOffloadedComponent_1_io_off_mem_req_bits_addr;
  wire[127:0] gTaggedDistributor_io_out_1_bits_data;
  wire[31:0] inputDist_io_out_1_bits_pageId;
  wire[31:0] gOffloadedComponent_io_off_mem_req_bits_addr;
  wire[127:0] gTaggedDistributor_io_out_0_bits_data;
  wire[31:0] inputDist_io_out_0_bits_pageId;
  wire gTaggedRRArbiter_io_out_valid;
  wire[31:0] inputDist_io_out_3_bits_pageId;
  wire[3:0] gOffloadedComponent_2_io_off_mem_req_bits_size;
  wire[3:0] gOffloadedComponent_1_io_off_mem_req_bits_size;
  wire[3:0] gOffloadedComponent_io_off_mem_req_bits_size;
  wire[127:0] gTaggedRRArbiter_io_out_bits_data;
  wire[127:0] gOffloadedComponent_3_io_off_mem_req_bits_data;
  wire[127:0] gOffloadedComponent_2_io_off_mem_req_bits_data;
  wire[127:0] gOffloadedComponent_1_io_off_mem_req_bits_data;
  wire[127:0] gOffloadedComponent_io_off_mem_req_bits_data;
  wire gTaggedRRArbiter_io_out_bits_cached;
  wire gOffloadedComponent_3_io_off_mem_req_bits_cached;
  wire gOffloadedComponent_2_io_off_mem_req_bits_cached;
  wire gOffloadedComponent_1_io_off_mem_req_bits_cached;
  wire gOffloadedComponent_io_off_mem_req_bits_cached;
  wire gTaggedRRArbiter_io_out_bits_rw;
  wire gOffloadedComponent_3_io_off_mem_req_bits_rw;
  wire gOffloadedComponent_2_io_off_mem_req_bits_rw;
  wire gOffloadedComponent_1_io_off_mem_req_bits_rw;
  wire gOffloadedComponent_io_off_mem_req_bits_rw;
  wire gTaggedDistributor_io_in_ready;
  wire gOffloadedComponent_3_io_off_mem_rep_ready;
  wire gOffloadedComponent_2_io_off_mem_rep_ready;
  wire gOffloadedComponent_1_io_off_mem_rep_ready;
  wire gOffloadedComponent_io_off_mem_rep_ready;
  wire[9:0] gTaggedRRArbiter_io_out_tag;
  wire[9:0] gOffloadedComponent_3_io_off_mem_req_tag;
  wire[9:0] gOffloadedComponent_2_io_off_mem_req_tag;
  wire[9:0] gOffloadedComponent_1_io_off_mem_req_tag;
  wire[9:0] gOffloadedComponent_io_off_mem_req_tag;
  wire[9:0] gTaggedRRArbiter_1_io_out_tag;
  wire[9:0] gOffloadedComponent_3_io_off_lock_req_tag;
  wire[9:0] gOffloadedComponent_2_io_off_lock_req_tag;
  wire[9:0] gOffloadedComponent_1_io_off_lock_req_tag;
  wire[9:0] gOffloadedComponent_io_off_lock_req_tag;
  wire gTaggedDistributor_1_io_out_3_valid;
  wire gTaggedRRArbiter_1_io_in_3_ready;
  wire gTaggedRRArbiter_io_in_3_ready;
  wire[9:0] outputArb_io_out_tag;
  wire[9:0] gOffloadedComponent_3_io_out_tag;
  wire[9:0] inputDist_io_out_3_tag;
  wire[9:0] gOffloadedComponent_2_io_out_tag;
  wire[9:0] inputDist_io_out_2_tag;
  wire[9:0] gOffloadedComponent_1_io_out_tag;
  wire[9:0] inputDist_io_out_1_tag;
  wire[9:0] gOffloadedComponent_io_out_tag;
  wire[9:0] inputDist_io_out_0_tag;
  wire outputArb_io_out_valid;
  wire[63:0] inputDist_io_out_0_bits_rankUpdate;
  wire[63:0] inputDist_io_out_1_bits_rankUpdate;
  wire[63:0] inputDist_io_out_2_bits_rankUpdate;
  wire[63:0] inputDist_io_out_3_bits_rankUpdate;

  assign io_in_ready = inputDist_io_in_ready;
  assign mainOff_lock_req_valid = gTaggedRRArbiter_1_io_out_valid;
  assign mainOff_mem_req_bits_size = gTaggedRRArbiter_io_out_bits_size;
  assign mainOff_lock_rep_ready = gTaggedDistributor_1_io_in_ready;
  assign mainOff_mem_req_bits_addr = gTaggedRRArbiter_io_out_bits_addr;
  assign mainOff_mem_req_valid = gTaggedRRArbiter_io_out_valid;
  assign mainOff_mem_req_bits_data = gTaggedRRArbiter_io_out_bits_data;
  assign mainOff_mem_req_bits_cached = gTaggedRRArbiter_io_out_bits_cached;
  assign mainOff_mem_req_bits_rw = gTaggedRRArbiter_io_out_bits_rw;
  assign mainOff_mem_rep_ready = gTaggedDistributor_io_in_ready;
  assign mainOff_mem_req_tag = gTaggedRRArbiter_io_out_tag;
  assign mainOff_lock_req_tag = gTaggedRRArbiter_1_io_out_tag;
  assign io_out_tag = outputArb_io_out_tag;
  assign io_out_valid = outputArb_io_out_valid;
  gOffloadedComponent_17 gOffloadedComponent(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_io_in_ready ),
       .io_in_valid( inputDist_io_out_0_valid ),
       .io_in_bits_done( inputDist_io_out_0_bits_done ),
       .io_in_bits_pageId( inputDist_io_out_0_bits_pageId ),
       .io_in_bits_rankUpdate( inputDist_io_out_0_bits_rankUpdate ),
       .io_in_tag( inputDist_io_out_0_tag ),
       .io_out_ready( outputArb_io_in_0_ready ),
       .io_out_valid( gOffloadedComponent_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( gOffloadedComponent_io_out_tag ),
       .pcIn0_valid(  ),
       .pcIn0_bits_request(  ),
       .pcIn0_bits_moduleId(  ),
       .pcIn0_bits_portId(  ),
       .pcIn0_bits_pcValue(  ),
       .pcIn0_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_0_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_0_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_0_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_0_tag ),
       .io_off_lock_req_ready( gTaggedRRArbiter_1_io_in_0_ready ),
       .io_off_lock_req_valid( gOffloadedComponent_io_off_lock_req_valid ),
       .io_off_lock_req_bits_id(  ),
       .io_off_lock_req_bits_op(  ),
       .io_off_lock_req_tag( gOffloadedComponent_io_off_lock_req_tag ),
       .io_off_lock_rep_ready( gOffloadedComponent_io_off_lock_rep_ready ),
       .io_off_lock_rep_valid( gTaggedDistributor_1_io_out_0_valid ),
       .io_off_lock_rep_bits_out(  ),
       .io_off_lock_rep_tag( gTaggedDistributor_1_io_out_0_tag ));
  gOffloadedComponent_18 gOffloadedComponent_1(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_1_io_in_ready ),
       .io_in_valid( inputDist_io_out_1_valid ),
       .io_in_bits_done( inputDist_io_out_1_bits_done ),
       .io_in_bits_pageId( inputDist_io_out_1_bits_pageId ),
       .io_in_bits_rankUpdate( inputDist_io_out_1_bits_rankUpdate ),
       .io_in_tag( inputDist_io_out_1_tag ),
       .io_out_ready( outputArb_io_in_1_ready ),
       .io_out_valid( gOffloadedComponent_1_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( gOffloadedComponent_1_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_1_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_1_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_1_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_1_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_1_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_1_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_1_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_1_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_1_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_1_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_1_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_1_tag ),
       .io_off_lock_req_ready( gTaggedRRArbiter_1_io_in_1_ready ),
       .io_off_lock_req_valid( gOffloadedComponent_1_io_off_lock_req_valid ),
       .io_off_lock_req_bits_id(  ),
       .io_off_lock_req_bits_op(  ),
       .io_off_lock_req_tag( gOffloadedComponent_1_io_off_lock_req_tag ),
       .io_off_lock_rep_ready( gOffloadedComponent_1_io_off_lock_rep_ready ),
       .io_off_lock_rep_valid( gTaggedDistributor_1_io_out_1_valid ),
       .io_off_lock_rep_bits_out(  ),
       .io_off_lock_rep_tag( gTaggedDistributor_1_io_out_1_tag ));
  gOffloadedComponent_19 gOffloadedComponent_2(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_2_io_in_ready ),
       .io_in_valid( inputDist_io_out_2_valid ),
       .io_in_bits_done( inputDist_io_out_2_bits_done ),
       .io_in_bits_pageId( inputDist_io_out_2_bits_pageId ),
       .io_in_bits_rankUpdate( inputDist_io_out_2_bits_rankUpdate ),
       .io_in_tag( inputDist_io_out_2_tag ),
       .io_out_ready( outputArb_io_in_2_ready ),
       .io_out_valid( gOffloadedComponent_2_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( gOffloadedComponent_2_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_2_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_2_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_2_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_2_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_2_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_2_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_2_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_2_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_2_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_2_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_2_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_2_tag ),
       .io_off_lock_req_ready( gTaggedRRArbiter_1_io_in_2_ready ),
       .io_off_lock_req_valid( gOffloadedComponent_2_io_off_lock_req_valid ),
       .io_off_lock_req_bits_id(  ),
       .io_off_lock_req_bits_op(  ),
       .io_off_lock_req_tag( gOffloadedComponent_2_io_off_lock_req_tag ),
       .io_off_lock_rep_ready( gOffloadedComponent_2_io_off_lock_rep_ready ),
       .io_off_lock_rep_valid( gTaggedDistributor_1_io_out_2_valid ),
       .io_off_lock_rep_bits_out(  ),
       .io_off_lock_rep_tag( gTaggedDistributor_1_io_out_2_tag ));
  gOffloadedComponent_20 gOffloadedComponent_3(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_3_io_in_ready ),
       .io_in_valid( inputDist_io_out_3_valid ),
       .io_in_bits_done( inputDist_io_out_3_bits_done ),
       .io_in_bits_pageId( inputDist_io_out_3_bits_pageId ),
       .io_in_bits_rankUpdate( inputDist_io_out_3_bits_rankUpdate ),
       .io_in_tag( inputDist_io_out_3_tag ),
       .io_out_ready( outputArb_io_in_3_ready ),
       .io_out_valid( gOffloadedComponent_3_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( gOffloadedComponent_3_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .pcOutN_valid(  ),
       .pcOutN_bits_request(  ),
       .pcOutN_bits_moduleId(  ),
       .pcOutN_bits_portId(  ),
       .pcOutN_bits_pcValue(  ),
       .pcOutN_bits_pcType(  ),
       .io_off_mem_req_ready( gTaggedRRArbiter_io_in_3_ready ),
       .io_off_mem_req_valid( gOffloadedComponent_3_io_off_mem_req_valid ),
       .io_off_mem_req_bits_addr( gOffloadedComponent_3_io_off_mem_req_bits_addr ),
       .io_off_mem_req_bits_rw( gOffloadedComponent_3_io_off_mem_req_bits_rw ),
       .io_off_mem_req_bits_cached( gOffloadedComponent_3_io_off_mem_req_bits_cached ),
       .io_off_mem_req_bits_data( gOffloadedComponent_3_io_off_mem_req_bits_data ),
       .io_off_mem_req_bits_size( gOffloadedComponent_3_io_off_mem_req_bits_size ),
       .io_off_mem_req_tag( gOffloadedComponent_3_io_off_mem_req_tag ),
       .io_off_mem_rep_ready( gOffloadedComponent_3_io_off_mem_rep_ready ),
       .io_off_mem_rep_valid( gTaggedDistributor_io_out_3_valid ),
       .io_off_mem_rep_bits_data( gTaggedDistributor_io_out_3_bits_data ),
       .io_off_mem_rep_tag( gTaggedDistributor_io_out_3_tag ),
       .io_off_lock_req_ready( gTaggedRRArbiter_1_io_in_3_ready ),
       .io_off_lock_req_valid( gOffloadedComponent_3_io_off_lock_req_valid ),
       .io_off_lock_req_bits_id(  ),
       .io_off_lock_req_bits_op(  ),
       .io_off_lock_req_tag( gOffloadedComponent_3_io_off_lock_req_tag ),
       .io_off_lock_rep_ready( gOffloadedComponent_3_io_off_lock_rep_ready ),
       .io_off_lock_rep_valid( gTaggedDistributor_1_io_out_3_valid ),
       .io_off_lock_rep_bits_out(  ),
       .io_off_lock_rep_tag( gTaggedDistributor_1_io_out_3_tag ));
  RRDistributorComponent_1 inputDist(.clk(clk), .reset(reset),
       .io_out_0_ready( gOffloadedComponent_io_in_ready ),
       .io_out_0_valid( inputDist_io_out_0_valid ),
       .io_out_0_bits_done( inputDist_io_out_0_bits_done ),
       .io_out_0_bits_pageId( inputDist_io_out_0_bits_pageId ),
       .io_out_0_bits_rankUpdate( inputDist_io_out_0_bits_rankUpdate ),
       .io_out_0_tag( inputDist_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_in_ready ),
       .io_out_1_valid( inputDist_io_out_1_valid ),
       .io_out_1_bits_done( inputDist_io_out_1_bits_done ),
       .io_out_1_bits_pageId( inputDist_io_out_1_bits_pageId ),
       .io_out_1_bits_rankUpdate( inputDist_io_out_1_bits_rankUpdate ),
       .io_out_1_tag( inputDist_io_out_1_tag ),
       .io_out_2_ready( gOffloadedComponent_2_io_in_ready ),
       .io_out_2_valid( inputDist_io_out_2_valid ),
       .io_out_2_bits_done( inputDist_io_out_2_bits_done ),
       .io_out_2_bits_pageId( inputDist_io_out_2_bits_pageId ),
       .io_out_2_bits_rankUpdate( inputDist_io_out_2_bits_rankUpdate ),
       .io_out_2_tag( inputDist_io_out_2_tag ),
       .io_out_3_ready( gOffloadedComponent_3_io_in_ready ),
       .io_out_3_valid( inputDist_io_out_3_valid ),
       .io_out_3_bits_done( inputDist_io_out_3_bits_done ),
       .io_out_3_bits_pageId( inputDist_io_out_3_bits_pageId ),
       .io_out_3_bits_rankUpdate( inputDist_io_out_3_bits_rankUpdate ),
       .io_out_3_tag( inputDist_io_out_3_tag ),
       .io_in_ready( inputDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
  RRAggregatorComponent_1 outputArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( outputArb_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( outputArb_io_out_tag ),
       .io_in_0_ready( outputArb_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_out_valid ),
       .io_in_0_bits_out(  ),
       .io_in_0_tag( gOffloadedComponent_io_out_tag ),
       .io_in_1_ready( outputArb_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_out_valid ),
       .io_in_1_bits_out(  ),
       .io_in_1_tag( gOffloadedComponent_1_io_out_tag ),
       .io_in_2_ready( outputArb_io_in_2_ready ),
       .io_in_2_valid( gOffloadedComponent_2_io_out_valid ),
       .io_in_2_bits_out(  ),
       .io_in_2_tag( gOffloadedComponent_2_io_out_tag ),
       .io_in_3_ready( outputArb_io_in_3_ready ),
       .io_in_3_valid( gOffloadedComponent_3_io_out_valid ),
       .io_in_3_bits_out(  ),
       .io_in_3_tag( gOffloadedComponent_3_io_out_tag ),
       .io_chosen(  ));
  gTaggedRRArbiter_1 gTaggedRRArbiter(.clk(clk), .reset(reset),
       .io_out_ready( mainOff_mem_req_ready ),
       .io_out_valid( gTaggedRRArbiter_io_out_valid ),
       .io_out_bits_addr( gTaggedRRArbiter_io_out_bits_addr ),
       .io_out_bits_rw( gTaggedRRArbiter_io_out_bits_rw ),
       .io_out_bits_cached( gTaggedRRArbiter_io_out_bits_cached ),
       .io_out_bits_data( gTaggedRRArbiter_io_out_bits_data ),
       .io_out_bits_size( gTaggedRRArbiter_io_out_bits_size ),
       .io_out_tag( gTaggedRRArbiter_io_out_tag ),
       .io_in_0_ready( gTaggedRRArbiter_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_off_mem_req_valid ),
       .io_in_0_bits_addr( gOffloadedComponent_io_off_mem_req_bits_addr ),
       .io_in_0_bits_rw( gOffloadedComponent_io_off_mem_req_bits_rw ),
       .io_in_0_bits_cached( gOffloadedComponent_io_off_mem_req_bits_cached ),
       .io_in_0_bits_data( gOffloadedComponent_io_off_mem_req_bits_data ),
       .io_in_0_bits_size( gOffloadedComponent_io_off_mem_req_bits_size ),
       .io_in_0_tag( gOffloadedComponent_io_off_mem_req_tag ),
       .io_in_1_ready( gTaggedRRArbiter_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_off_mem_req_valid ),
       .io_in_1_bits_addr( gOffloadedComponent_1_io_off_mem_req_bits_addr ),
       .io_in_1_bits_rw( gOffloadedComponent_1_io_off_mem_req_bits_rw ),
       .io_in_1_bits_cached( gOffloadedComponent_1_io_off_mem_req_bits_cached ),
       .io_in_1_bits_data( gOffloadedComponent_1_io_off_mem_req_bits_data ),
       .io_in_1_bits_size( gOffloadedComponent_1_io_off_mem_req_bits_size ),
       .io_in_1_tag( gOffloadedComponent_1_io_off_mem_req_tag ),
       .io_in_2_ready( gTaggedRRArbiter_io_in_2_ready ),
       .io_in_2_valid( gOffloadedComponent_2_io_off_mem_req_valid ),
       .io_in_2_bits_addr( gOffloadedComponent_2_io_off_mem_req_bits_addr ),
       .io_in_2_bits_rw( gOffloadedComponent_2_io_off_mem_req_bits_rw ),
       .io_in_2_bits_cached( gOffloadedComponent_2_io_off_mem_req_bits_cached ),
       .io_in_2_bits_data( gOffloadedComponent_2_io_off_mem_req_bits_data ),
       .io_in_2_bits_size( gOffloadedComponent_2_io_off_mem_req_bits_size ),
       .io_in_2_tag( gOffloadedComponent_2_io_off_mem_req_tag ),
       .io_in_3_ready( gTaggedRRArbiter_io_in_3_ready ),
       .io_in_3_valid( gOffloadedComponent_3_io_off_mem_req_valid ),
       .io_in_3_bits_addr( gOffloadedComponent_3_io_off_mem_req_bits_addr ),
       .io_in_3_bits_rw( gOffloadedComponent_3_io_off_mem_req_bits_rw ),
       .io_in_3_bits_cached( gOffloadedComponent_3_io_off_mem_req_bits_cached ),
       .io_in_3_bits_data( gOffloadedComponent_3_io_off_mem_req_bits_data ),
       .io_in_3_bits_size( gOffloadedComponent_3_io_off_mem_req_bits_size ),
       .io_in_3_tag( gOffloadedComponent_3_io_off_mem_req_tag ),
       .io_chosen(  ));
  gTaggedRRArbiter_2 gTaggedRRArbiter_1(.clk(clk), .reset(reset),
       .io_out_ready( mainOff_lock_req_ready ),
       .io_out_valid( gTaggedRRArbiter_1_io_out_valid ),
       .io_out_bits_id(  ),
       .io_out_bits_op(  ),
       .io_out_tag( gTaggedRRArbiter_1_io_out_tag ),
       .io_in_0_ready( gTaggedRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_off_lock_req_valid ),
       .io_in_0_bits_id(  ),
       .io_in_0_bits_op(  ),
       .io_in_0_tag( gOffloadedComponent_io_off_lock_req_tag ),
       .io_in_1_ready( gTaggedRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_off_lock_req_valid ),
       .io_in_1_bits_id(  ),
       .io_in_1_bits_op(  ),
       .io_in_1_tag( gOffloadedComponent_1_io_off_lock_req_tag ),
       .io_in_2_ready( gTaggedRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( gOffloadedComponent_2_io_off_lock_req_valid ),
       .io_in_2_bits_id(  ),
       .io_in_2_bits_op(  ),
       .io_in_2_tag( gOffloadedComponent_2_io_off_lock_req_tag ),
       .io_in_3_ready( gTaggedRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( gOffloadedComponent_3_io_off_lock_req_valid ),
       .io_in_3_bits_id(  ),
       .io_in_3_bits_op(  ),
       .io_in_3_tag( gOffloadedComponent_3_io_off_lock_req_tag ),
       .io_chosen(  ));
  gTaggedDistributor_1 gTaggedDistributor(
       .io_out_0_ready( gOffloadedComponent_io_off_mem_rep_ready ),
       .io_out_0_valid( gTaggedDistributor_io_out_0_valid ),
       .io_out_0_bits_data( gTaggedDistributor_io_out_0_bits_data ),
       .io_out_0_tag( gTaggedDistributor_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_off_mem_rep_ready ),
       .io_out_1_valid( gTaggedDistributor_io_out_1_valid ),
       .io_out_1_bits_data( gTaggedDistributor_io_out_1_bits_data ),
       .io_out_1_tag( gTaggedDistributor_io_out_1_tag ),
       .io_out_2_ready( gOffloadedComponent_2_io_off_mem_rep_ready ),
       .io_out_2_valid( gTaggedDistributor_io_out_2_valid ),
       .io_out_2_bits_data( gTaggedDistributor_io_out_2_bits_data ),
       .io_out_2_tag( gTaggedDistributor_io_out_2_tag ),
       .io_out_3_ready( gOffloadedComponent_3_io_off_mem_rep_ready ),
       .io_out_3_valid( gTaggedDistributor_io_out_3_valid ),
       .io_out_3_bits_data( gTaggedDistributor_io_out_3_bits_data ),
       .io_out_3_tag( gTaggedDistributor_io_out_3_tag ),
       .io_in_ready( gTaggedDistributor_io_in_ready ),
       .io_in_valid( mainOff_mem_rep_valid ),
       .io_in_bits_data( mainOff_mem_rep_bits_data ),
       .io_in_tag( mainOff_mem_rep_tag ),
       .io_chosen(  ));
  gTaggedDistributor_2 gTaggedDistributor_1(
       .io_out_0_ready( gOffloadedComponent_io_off_lock_rep_ready ),
       .io_out_0_valid( gTaggedDistributor_1_io_out_0_valid ),
       .io_out_0_bits_out(  ),
       .io_out_0_tag( gTaggedDistributor_1_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_off_lock_rep_ready ),
       .io_out_1_valid( gTaggedDistributor_1_io_out_1_valid ),
       .io_out_1_bits_out(  ),
       .io_out_1_tag( gTaggedDistributor_1_io_out_1_tag ),
       .io_out_2_ready( gOffloadedComponent_2_io_off_lock_rep_ready ),
       .io_out_2_valid( gTaggedDistributor_1_io_out_2_valid ),
       .io_out_2_bits_out(  ),
       .io_out_2_tag( gTaggedDistributor_1_io_out_2_tag ),
       .io_out_3_ready( gOffloadedComponent_3_io_off_lock_rep_ready ),
       .io_out_3_valid( gTaggedDistributor_1_io_out_3_valid ),
       .io_out_3_bits_out(  ),
       .io_out_3_tag( gTaggedDistributor_1_io_out_3_tag ),
       .io_in_ready( gTaggedDistributor_1_io_in_ready ),
       .io_in_valid( mainOff_lock_rep_valid ),
       .io_in_bits_out(  ),
       .io_in_tag( mainOff_lock_rep_tag ),
       .io_chosen(  ));
endmodule

module lockModel(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_id,
    input  io_in_bits_op,
    input [9:0] io_in_tag,
    input  outputReg_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] outputReg_tag;
  wire T0;
  wire T1;
  reg[0:0] outputReg_valid;
  wire T2;
  wire[9:0] T3;
  wire[9:0] T4;

  assign io_out_tag = outputReg_tag;
  assign T0 = outputReg_ready || T1;
  assign T1 = ! outputReg_valid;
  assign T2 = T0 ? io_in_valid : outputReg_valid;
  assign io_out_valid = outputReg_valid;
  assign io_in_ready = outputReg_ready;
  assign T4 = T0 ? io_in_tag : outputReg_tag;

  always @(posedge clk) begin
    if(reset) begin
      outputReg_tag <= T3;
    end else if(T0) begin
      outputReg_tag <= T4;
    end
    if(reset) begin
      outputReg_valid <= 1'h0/* 0*/;
    end else if(T0) begin
      outputReg_valid <= T2;
    end
  end
endmodule

module gOffloadedComponent_21(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_mem_req_ready,
    output mainOff_mem_req_valid,
    output[31:0] mainOff_mem_req_bits_addr,
    output mainOff_mem_req_bits_rw,
    output mainOff_mem_req_bits_cached,
    output[127:0] mainOff_mem_req_bits_data,
    output[3:0] mainOff_mem_req_bits_size,
    output[9:0] mainOff_mem_req_tag,
    output mainOff_mem_rep_ready,
    input  mainOff_mem_rep_valid,
    input [127:0] mainOff_mem_rep_bits_data,
    input [9:0] mainOff_mem_rep_tag);

  wire mainComp_io_in_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_lock_req_valid;
  wire offComp_io_out_valid;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_lock_rep_ready;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire mainComp_mainOff_mem_req_valid;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_mainOff_lock_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_mem_req_bits_size = mainComp_mainOff_mem_req_bits_size;
  assign mainOff_mem_req_bits_addr = mainComp_mainOff_mem_req_bits_addr;
  assign mainOff_mem_req_valid = mainComp_mainOff_mem_req_valid;
  assign mainOff_mem_req_bits_data = mainComp_mainOff_mem_req_bits_data;
  assign mainOff_mem_req_bits_cached = mainComp_mainOff_mem_req_bits_cached;
  assign mainOff_mem_req_bits_rw = mainComp_mainOff_mem_req_bits_rw;
  assign mainOff_mem_rep_ready = mainComp_mainOff_mem_rep_ready;
  assign mainOff_mem_req_tag = mainComp_mainOff_mem_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gReplicatedComponent_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( mainOff_mem_req_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( mainOff_mem_rep_valid ),
       .mainOff_mem_rep_bits_data( mainOff_mem_rep_bits_data ),
       .mainOff_mem_rep_tag( mainOff_mem_rep_tag ),
       .mainOff_lock_req_ready( offComp_io_in_ready ),
       .mainOff_lock_req_valid( mainComp_mainOff_lock_req_valid ),
       .mainOff_lock_req_bits_id(  ),
       .mainOff_lock_req_bits_op(  ),
       .mainOff_lock_req_tag( mainComp_mainOff_lock_req_tag ),
       .mainOff_lock_rep_ready( mainComp_mainOff_lock_rep_ready ),
       .mainOff_lock_rep_valid( offComp_io_out_valid ),
       .mainOff_lock_rep_bits_out(  ),
       .mainOff_lock_rep_tag( offComp_io_out_tag ));
  lockModel offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_lock_req_valid ),
       .io_in_bits_id(  ),
       .io_in_bits_op(  ),
       .io_in_tag( mainComp_mainOff_lock_req_tag ),
       .outputReg_ready( mainComp_mainOff_lock_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_56(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_57(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_58(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module cache_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_cacheMissPipe_req_ready,
    output mainOff_cacheMissPipe_req_valid,
    output[31:0] mainOff_cacheMissPipe_req_bits,
    output[9:0] mainOff_cacheMissPipe_req_tag,
    output mainOff_cacheMissPipe_rep_ready,
    input  mainOff_cacheMissPipe_rep_valid,
    input [31:0] mainOff_cacheMissPipe_rep_bits,
    input [9:0] mainOff_cacheMissPipe_rep_tag,
    input  mainOff_dram_req_ready,
    output mainOff_dram_req_valid,
    output[31:0] mainOff_dram_req_bits_addr,
    output mainOff_dram_req_bits_rw,
    output mainOff_dram_req_bits_cached,
    output[127:0] mainOff_dram_req_bits_data,
    output[3:0] mainOff_dram_req_bits_size,
    output[9:0] mainOff_dram_req_tag,
    output mainOff_dram_rep_ready,
    input  mainOff_dram_rep_valid,
    input [127:0] mainOff_dram_rep_bits_data,
    input [9:0] mainOff_dram_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire[9:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T6;
  reg[0:0] subStateTh_2;
  wire T7;
  wire T8;
  wire T9;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T10;
  wire AllOffloadsValid_2;
  wire T11;
  wire T12;
  wire T13;
  reg[0:0] dramPortHadValidRequest_2;
  wire T14;
  wire T15;
  wire T16;
  wire dramPort_req_valid;
  wire T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire[7:0] T23;
  reg[7:0] State_2;
  wire T24;
  wire T25;
  wire T26;
  wire[2:0] T27;
  wire[5:0] T28;
  wire T29;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire T38;
  reg[7:0] State_1;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[7:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[31:0] T59;
  wire T60;
  wire T61;
  reg[0:0] inputReg_2_rw;
  wire T62;
  wire T63;
  wire[2:0] T64;
  wire[5:0] T65;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  reg[0:0] subStateTh_1;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire[1:0] T82;
  wire AllOffloadsReady;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] dramPortHadReadyRequest;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  reg[0:0] dram_ready_received;
  wire T92;
  wire T93;
  wire dramPort_req_ready;
  wire[31:0] dramPort_req_bits_addr;
  wire[31:0] T94;
  wire[165:0] T95;
  wire[165:0] T96;
  wire[165:0] T97;
  wire[3:0] T98;
  wire[3:0] T99;
  wire[3:0] T100;
  reg[3:0] inputReg_2_size;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire[127:0] T106;
  wire[127:0] T107;
  wire[127:0] T108;
  reg[127:0] outputReg_2_data;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire[55:0] T114;
  wire[31:0] T115;
  wire[31:0] T116;
  wire[31:0] T117;
  reg[31:0] inputReg_2_addr;
  wire[31:0] T118;
  wire[31:0] T119;
  wire[31:0] T120;
  wire[31:0] T121;
  reg[31:0] inputReg_1_addr;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[31:0] T126;
  wire[31:0] T127;
  wire[31:0] T128;
  wire T129;
  reg[31:0] inputReg_0_addr;
  wire T130;
  wire T131;
  wire[31:0] T132;
  wire T133;
  wire T134;
  wire[7:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire[31:0] T142;
  wire[31:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire[127:0] T147;
  wire[127:0] T148;
  wire[127:0] T149;
  wire[127:0] T150;
  wire[127:0] T151;
  wire[60:0] T152;
  wire[55:0] T153;
  wire[55:0] T154;
  wire[31:0] T155;
  wire[31:0] T156;
  wire[31:0] T157;
  reg[31:0] random_2;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  reg[31:0] burst_2;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire T175;
  wire[31:0] T176;
  wire[31:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  reg[31:0] burst_1;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[31:0] T184;
  wire[31:0] T185;
  wire T186;
  wire[31:0] T187;
  wire[31:0] T188;
  reg[31:0] burst_0;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire[31:0] T193;
  wire[31:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire[31:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[31:0] T205;
  wire[31:0] T206;
  wire T207;
  wire[31:0] T208;
  wire[31:0] T209;
  wire[31:0] T210;
  wire[31:0] T211;
  reg[31:0] random_1;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire T218;
  wire[31:0] T219;
  wire[31:0] T220;
  reg[31:0] random_0;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[31:0] T225;
  wire[31:0] T226;
  wire T227;
  wire[127:0] T228;
  wire[31:0] T229;
  wire[127:0] T230;
  wire[127:0] T231;
  wire[127:0] T232;
  wire T233;
  reg[127:0] outputReg_1_data;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire[127:0] T239;
  wire[127:0] T240;
  wire[127:0] T241;
  wire[127:0] T242;
  wire[127:0] T243;
  wire[127:0] T244;
  wire[127:0] T245;
  wire[127:0] T246;
  wire T247;
  reg[127:0] outputReg_0_data;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire[127:0] T253;
  wire[127:0] T254;
  wire[127:0] T255;
  wire[127:0] T256;
  wire[127:0] T257;
  wire[127:0] T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  reg[3:0] inputReg_1_size;
  wire[3:0] T262;
  wire[3:0] T263;
  wire[3:0] T264;
  reg[3:0] inputReg_0_size;
  wire[3:0] T265;
  wire[127:0] T266;
  wire[127:0] T267;
  wire[127:0] T268;
  reg[127:0] inputReg_2_data;
  wire[127:0] T269;
  wire[127:0] T270;
  wire[127:0] T271;
  wire[127:0] T272;
  reg[127:0] inputReg_1_data;
  wire[127:0] T273;
  wire[127:0] T274;
  wire[127:0] T275;
  reg[127:0] inputReg_0_data;
  wire[127:0] T276;
  wire T277;
  wire T278;
  reg[0:0] inputReg_2_cached;
  wire T279;
  wire T280;
  wire T281;
  reg[0:0] inputReg_1_cached;
  wire T282;
  wire T283;
  reg[0:0] inputReg_0_cached;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  reg[0:0] inputReg_1_rw;
  wire T289;
  wire T290;
  reg[0:0] inputReg_0_rw;
  wire T291;
  wire[31:0] T292;
  wire[31:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[31:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire T300;
  wire T301;
  wire[7:0] T302;
  wire T303;
  wire dramPort_rep_ready;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire cacheMissPipePort_req_valid;
  wire T308;
  wire T309;
  wire T310;
  wire[7:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  reg[0:0] cacheMissPipe_valid_received_2;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[9:0] T321;
  wire[9:0] cacheMissPipePort_rep_tag;
  wire cacheMissPipePort_rep_ready;
  wire[9:0] cacheMissPipePort_req_tag;
  wire[9:0] T322;
  wire cacheMissPipePort_rep_valid;
  wire T323;
  wire T324;
  wire[4:0] T325;
  wire T326;
  wire T327;
  reg[0:0] cacheMissPipe_valid_received_1;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[9:0] T332;
  wire T333;
  wire T334;
  wire[4:0] T335;
  wire T336;
  reg[0:0] cacheMissPipe_valid_received_0;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire[9:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  reg[0:0] cacheMissPipePortHadReadyRequest;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  reg[0:0] cacheMissPipe_ready_received;
  wire T351;
  wire T352;
  wire cacheMissPipePort_req_ready;
  wire T353;
  wire T354;
  wire T355;
  reg[7:0] State_0;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire[7:0] T373;
  wire[7:0] T374;
  wire[7:0] T375;
  wire[7:0] T376;
  wire[7:0] T377;
  wire[7:0] T378;
  wire[7:0] T379;
  wire[7:0] T380;
  wire[7:0] T381;
  wire[7:0] T382;
  wire[7:0] T383;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[7:0] T386;
  wire[7:0] T387;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T388;
  wire[7:0] T389;
  wire[7:0] T390;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T391;
  wire[7:0] T392;
  wire[7:0] T393;
  wire[7:0] T394;
  wire[7:0] T395;
  wire T396;
  reg[0:0] subStateTh_0;
  wire T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire[1:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire[31:0] T414;
  wire[31:0] T415;
  wire[31:0] T416;
  reg[31:0] cachedAddr_2;
  wire T417;
  wire T418;
  wire[31:0] T419;
  wire[31:0] T420;
  wire[31:0] ct;
  wire[31:0] T421;
  wire[31:0] T422;
  wire[31:0] T423;
  reg[31:0] cachedAddr_1;
  wire T424;
  wire[31:0] T425;
  wire[31:0] T426;
  wire[31:0] T427;
  wire[31:0] T428;
  reg[31:0] cachedAddr_0;
  wire T429;
  wire[31:0] T430;
  wire[31:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[7:0] T436;
  wire[7:0] T437;
  wire[7:0] T438;
  wire[7:0] T439;
  wire[7:0] T440;
  wire[7:0] T441;
  wire[7:0] T442;
  wire[7:0] T443;
  wire[7:0] T444;
  wire[7:0] T445;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T448;
  wire[7:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  reg[0:0] dram_valid_received_2;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[9:0] T486;
  wire[9:0] dramPort_rep_tag;
  wire[9:0] dramPort_req_tag;
  wire[9:0] T487;
  wire dramPort_rep_valid;
  wire T488;
  wire T489;
  wire[4:0] T490;
  wire T491;
  wire T492;
  reg[0:0] dram_valid_received_1;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire[9:0] T497;
  wire T498;
  wire T499;
  wire[4:0] T500;
  wire T501;
  reg[0:0] dram_valid_received_0;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire[9:0] T506;
  wire T507;
  wire T508;
  wire[4:0] T509;
  wire T510;
  wire T511;
  wire[4:0] T512;
  wire T513;
  wire T514;
  wire[4:0] T515;
  wire T516;
  wire T517;
  wire T518;
  wire[9:0] T519;
  wire T520;
  wire T521;
  reg[0:0] cacheMissPipePortHadValidRequest_2;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[4:0] T526;
  wire T527;
  wire T528;
  wire[4:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire[9:0] T533;
  wire T534;
  wire T535;
  wire AllOffloadsValid_1;
  wire T536;
  wire T537;
  wire T538;
  reg[0:0] dramPortHadValidRequest_1;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire[4:0] T543;
  wire T544;
  wire T545;
  wire[4:0] T546;
  wire T547;
  wire T548;
  wire T549;
  wire[9:0] T550;
  wire T551;
  wire T552;
  reg[0:0] cacheMissPipePortHadValidRequest_1;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire[4:0] T557;
  wire T558;
  wire T559;
  wire[4:0] T560;
  wire T561;
  wire T562;
  wire T563;
  wire[9:0] T564;
  wire T565;
  wire T566;
  wire AllOffloadsValid_0;
  wire T567;
  wire T568;
  wire T569;
  reg[0:0] dramPortHadValidRequest_0;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[4:0] T574;
  wire T575;
  wire T576;
  wire[4:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire[9:0] T581;
  wire T582;
  wire T583;
  reg[0:0] cacheMissPipePortHadValidRequest_0;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[4:0] T588;
  wire T589;
  wire T590;
  wire[4:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[9:0] T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[9:0] inputTag_2;
  wire[9:0] T607;
  wire[9:0] T608;
  wire[9:0] T609;
  wire[9:0] T610;
  reg[9:0] inputTag_1;
  wire[9:0] T611;
  wire[9:0] T612;
  wire[9:0] T613;
  reg[9:0] inputTag_0;
  wire[9:0] T614;

  assign io_out_tag = T0;
  assign T0 = T608 | T1;
  assign T1 = inputTag_2 & T2;
  assign T2 = {4'ha/* 10*/{T3}};
  assign T3 = T4[2'h2/* 2*/];
  assign T4 = T5[2'h2/* 2*/:1'h0/* 0*/];
  assign T5 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T6 = subStateTh_2 == 1'h0/* 0*/;
  assign T7 = T598 ? 1'h1/* 1*/ : T8;
  assign T8 = T9 ? 1'h0/* 0*/ : subStateTh_2;
  assign T9 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T10 = T534 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T11;
  assign T11 = T520 && T12;
  assign T12 = T516 || T13;
  assign T13 = ! dramPortHadValidRequest_2;
  assign T14 = T513 && T15;
  assign T15 = dramPortHadValidRequest_2 || T16;
  assign T16 = T511 && dramPort_req_valid;
  assign dramPort_req_valid = T17;
  assign T17 = T478 && T18;
  assign T18 = T477 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = T472 | T22;
  assign T22 = State_2 & T23;
  assign T23 = {4'h8/* 8*/{T3}};
  assign T24 = T451 || T25;
  assign T25 = T29 && T26;
  assign T26 = T27[2'h2/* 2*/];
  assign T27 = T28[2'h2/* 2*/:1'h0/* 0*/];
  assign T28 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T29 = T450 && T30;
  assign T30 = T32 == T31;
  assign T31 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T32 = T35 | T33;
  assign T33 = State_2 & T34;
  assign T34 = {4'h8/* 8*/{T26}};
  assign T35 = T448 | T36;
  assign T36 = State_1 & T37;
  assign T37 = {4'h8/* 8*/{T38}};
  assign T38 = T27[1'h1/* 1*/];
  assign T39 = T41 || T40;
  assign T40 = T29 && T38;
  assign T41 = T47 || T42;
  assign T42 = T43 && T38;
  assign T43 = T46 && T44;
  assign T44 = T32 == T45;
  assign T45 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T46 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T47 = T53 || T48;
  assign T48 = T49 && T38;
  assign T49 = T52 && T50;
  assign T50 = T32 == T51;
  assign T51 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T52 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T53 = T432 || T54;
  assign T54 = T55 && T38;
  assign T55 = T133 && T56;
  assign T56 = ! T57;
  assign T57 = T413 || T58;
  assign T58 = T59 == 32'h1/* 1*/;
  assign T59 = {31'h0/* 0*/, T60};
  assign T60 = T410 | T61;
  assign T61 = inputReg_2_rw & T26;
  assign T62 = T124 && T63;
  assign T63 = T64[2'h2/* 2*/];
  assign T64 = T65[2'h2/* 2*/:1'h0/* 0*/];
  assign T65 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T66 = T68 && T67;
  assign T67 = State_2 == 8'h0/* 0*/;
  assign T68 = subStateTh_2 == 1'h0/* 0*/;
  assign T69 = T71 && T70;
  assign T70 = State_1 == 8'h0/* 0*/;
  assign T71 = subStateTh_1 == 1'h0/* 0*/;
  assign T72 = T76 ? 1'h1/* 1*/ : T73;
  assign T73 = T74 ? 1'h0/* 0*/ : subStateTh_1;
  assign T74 = T75 == vThreadEncoder_io_chosen;
  assign T75 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T76 = T78 && T77;
  assign T77 = State_1 != 8'hff/* 255*/;
  assign T78 = T80 && T79;
  assign T79 = State_1 != 8'h0/* 0*/;
  assign T80 = AllOffloadsReady && T81;
  assign T81 = T82 == rThreadEncoder_io_chosen;
  assign T82 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign AllOffloadsReady = T83;
  assign T83 = T305 && T84;
  assign T84 = T91 || T85;
  assign T85 = T87 && T86;
  assign T86 = ! dramPort_req_valid;
  assign T87 = ! dramPortHadReadyRequest;
  assign T88 = T90 && T89;
  assign T89 = dramPortHadReadyRequest || dramPort_req_valid;
  assign T90 = ! AllOffloadsReady;
  assign T91 = dramPort_req_ready || dram_ready_received;
  assign T92 = T304 && T93;
  assign T93 = dram_ready_received || dramPort_req_ready;
  assign dramPort_req_ready = mainOff_dram_req_ready;
  assign mainOff_dram_req_valid = dramPort_req_valid;
  assign mainOff_dram_req_bits_addr = dramPort_req_bits_addr;
  assign dramPort_req_bits_addr = T94;
  assign T94 = T95[8'ha5/* 165*/:8'h86/* 134*/];
  assign T95 = T300 ? T97 : T96;
  assign T96 = {134'h0/* 0*/, 32'h0/* 0*/};
  assign T97 = {T292, T285, T277, T266, T98};
  assign T98 = T259 | T99;
  assign T99 = inputReg_2_size & T100;
  assign T100 = {3'h4/* 4*/{T3}};
  assign T101 = T62 ? io_in_bits_size : inputReg_2_size;
  assign io_out_valid = T102;
  assign T102 = T104 && T103;
  assign T103 = T21 == 8'hff/* 255*/;
  assign T104 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_in_ready = T105;
  assign T105 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_data = T106;
  assign T106 = T230 | T107;
  assign T107 = outputReg_2_data & T108;
  assign T108 = {8'h80/* 128*/{T3}};
  assign T109 = T137 || T110;
  assign T110 = T111 && T26;
  assign T111 = T133 && T112;
  assign T112 = ! T113;
  assign T113 = T114 <= 56'h1000000/* 16777216*/;
  assign T114 = {24'h0/* 0*/, T115};
  assign T115 = T119 | T116;
  assign T116 = inputReg_2_addr & T117;
  assign T117 = {6'h20/* 32*/{T26}};
  assign T118 = T62 ? io_in_bits_addr : inputReg_2_addr;
  assign T119 = T127 | T120;
  assign T120 = inputReg_1_addr & T121;
  assign T121 = {6'h20/* 32*/{T38}};
  assign T122 = T124 && T123;
  assign T123 = T64[1'h1/* 1*/];
  assign T124 = T125 && io_in_valid;
  assign T125 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T126 = T122 ? io_in_bits_addr : inputReg_1_addr;
  assign T127 = inputReg_0_addr & T128;
  assign T128 = {6'h20/* 32*/{T129}};
  assign T129 = T27[1'h0/* 0*/];
  assign T130 = T124 && T131;
  assign T131 = T64[1'h0/* 0*/];
  assign T132 = T130 ? io_in_bits_addr : inputReg_0_addr;
  assign T133 = T136 && T134;
  assign T134 = T32 == T135;
  assign T135 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T136 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T137 = T145 || T138;
  assign T138 = T139 && T26;
  assign T139 = T144 && T140;
  assign T140 = ! T141;
  assign T141 = T142 == 32'h0/* 0*/;
  assign T142 = T143 & 32'h1/* 1*/;
  assign T143 = T115 >> 32'h2/* 2*/;
  assign T144 = T133 && T113;
  assign T145 = T146 && T26;
  assign T146 = T144 && T141;
  assign T147 = T110 ? T228 : T148;
  assign T148 = T138 ? T151 : T149;
  assign T149 = T145 ? T150 : outputReg_2_data;
  assign T150 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T151 = {67'h0/* 0*/, T152};
  assign T152 = T153 << 32'h5/* 5*/;
  assign T153 = 56'h1000000/* 16777216*/ + T154;
  assign T154 = {24'h0/* 0*/, T155};
  assign T155 = T209 | T156;
  assign T156 = random_2 & T157;
  assign T157 = {6'h20/* 32*/{T26}};
  assign T158 = T200 || T159;
  assign T159 = T160 && T26;
  assign T160 = T196 && T161;
  assign T161 = T162 == 32'h1/* 1*/;
  assign T162 = T177 | T163;
  assign T163 = burst_2 & T164;
  assign T164 = {6'h20/* 32*/{T26}};
  assign T165 = T170 || T166;
  assign T166 = T167 && T26;
  assign T167 = T146 && T168;
  assign T168 = ! T169;
  assign T169 = T162 == 32'h1/* 1*/;
  assign T170 = T62 || T171;
  assign T171 = T172 && T26;
  assign T172 = T146 && T169;
  assign T173 = T166 ? T176 : T174;
  assign T174 = T175 ? 32'h1/* 1*/ : burst_2;
  assign T175 = T62 || T171;
  assign T176 = T162 + 32'h1/* 1*/;
  assign T177 = T187 | T178;
  assign T178 = burst_1 & T179;
  assign T179 = {6'h20/* 32*/{T38}};
  assign T180 = T182 || T181;
  assign T181 = T167 && T38;
  assign T182 = T122 || T183;
  assign T183 = T172 && T38;
  assign T184 = T181 ? T176 : T185;
  assign T185 = T186 ? 32'h1/* 1*/ : burst_1;
  assign T186 = T122 || T183;
  assign T187 = burst_0 & T188;
  assign T188 = {6'h20/* 32*/{T129}};
  assign T189 = T191 || T190;
  assign T190 = T167 && T129;
  assign T191 = T130 || T192;
  assign T192 = T172 && T129;
  assign T193 = T190 ? T176 : T194;
  assign T194 = T195 ? 32'h1/* 1*/ : burst_0;
  assign T195 = T130 || T192;
  assign T196 = T146 && T197;
  assign T197 = ! T198;
  assign T198 = T155 == T199;
  assign T199 = {1'h0/* 0*/, 31'h2/* 2*/};
  assign T200 = T62 || T201;
  assign T201 = T202 && T26;
  assign T202 = T204 && T203;
  assign T203 = T162 == 32'h1/* 1*/;
  assign T204 = T146 && T198;
  assign T205 = T159 ? T208 : T206;
  assign T206 = T207 ? 32'h1/* 1*/ : random_2;
  assign T207 = T62 || T201;
  assign T208 = T155 + 32'h1/* 1*/;
  assign T209 = T219 | T210;
  assign T210 = random_1 & T211;
  assign T211 = {6'h20/* 32*/{T38}};
  assign T212 = T214 || T213;
  assign T213 = T160 && T38;
  assign T214 = T122 || T215;
  assign T215 = T202 && T38;
  assign T216 = T213 ? T208 : T217;
  assign T217 = T218 ? 32'h1/* 1*/ : random_1;
  assign T218 = T122 || T215;
  assign T219 = random_0 & T220;
  assign T220 = {6'h20/* 32*/{T129}};
  assign T221 = T223 || T222;
  assign T222 = T160 && T129;
  assign T223 = T130 || T224;
  assign T224 = T202 && T129;
  assign T225 = T222 ? T208 : T226;
  assign T226 = T227 ? 32'h1/* 1*/ : random_0;
  assign T227 = T130 || T224;
  assign T228 = {96'h0/* 0*/, T229};
  assign T229 = T115 + 32'h3e8/* 1000*/;
  assign T230 = T245 | T231;
  assign T231 = outputReg_1_data & T232;
  assign T232 = {8'h80/* 128*/{T233}};
  assign T233 = T4[1'h1/* 1*/];
  assign T234 = T236 || T235;
  assign T235 = T111 && T38;
  assign T236 = T238 || T237;
  assign T237 = T139 && T38;
  assign T238 = T146 && T38;
  assign T239 = T235 ? T244 : T240;
  assign T240 = T237 ? T243 : T241;
  assign T241 = T238 ? T242 : outputReg_1_data;
  assign T242 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T243 = {67'h0/* 0*/, T152};
  assign T244 = {96'h0/* 0*/, T229};
  assign T245 = outputReg_0_data & T246;
  assign T246 = {8'h80/* 128*/{T247}};
  assign T247 = T4[1'h0/* 0*/];
  assign T248 = T250 || T249;
  assign T249 = T111 && T129;
  assign T250 = T252 || T251;
  assign T251 = T139 && T129;
  assign T252 = T146 && T129;
  assign T253 = T249 ? T258 : T254;
  assign T254 = T251 ? T257 : T255;
  assign T255 = T252 ? T256 : outputReg_0_data;
  assign T256 = {96'h0/* 0*/, 32'h5/* 5*/};
  assign T257 = {67'h0/* 0*/, T152};
  assign T258 = {96'h0/* 0*/, T229};
  assign T259 = T263 | T260;
  assign T260 = inputReg_1_size & T261;
  assign T261 = {3'h4/* 4*/{T233}};
  assign T262 = T122 ? io_in_bits_size : inputReg_1_size;
  assign T263 = inputReg_0_size & T264;
  assign T264 = {3'h4/* 4*/{T247}};
  assign T265 = T130 ? io_in_bits_size : inputReg_0_size;
  assign T266 = T270 | T267;
  assign T267 = inputReg_2_data & T268;
  assign T268 = {8'h80/* 128*/{T3}};
  assign T269 = T62 ? io_in_bits_data : inputReg_2_data;
  assign T270 = T274 | T271;
  assign T271 = inputReg_1_data & T272;
  assign T272 = {8'h80/* 128*/{T233}};
  assign T273 = T122 ? io_in_bits_data : inputReg_1_data;
  assign T274 = inputReg_0_data & T275;
  assign T275 = {8'h80/* 128*/{T247}};
  assign T276 = T130 ? io_in_bits_data : inputReg_0_data;
  assign T277 = T280 | T278;
  assign T278 = inputReg_2_cached & T3;
  assign T279 = T62 ? io_in_bits_cached : inputReg_2_cached;
  assign T280 = T283 | T281;
  assign T281 = inputReg_1_cached & T233;
  assign T282 = T122 ? io_in_bits_cached : inputReg_1_cached;
  assign T283 = inputReg_0_cached & T247;
  assign T284 = T130 ? io_in_bits_cached : inputReg_0_cached;
  assign T285 = T287 | T286;
  assign T286 = inputReg_2_rw & T3;
  assign T287 = T290 | T288;
  assign T288 = inputReg_1_rw & T233;
  assign T289 = T122 ? io_in_bits_rw : inputReg_1_rw;
  assign T290 = inputReg_0_rw & T247;
  assign T291 = T130 ? io_in_bits_rw : inputReg_0_rw;
  assign T292 = T295 | T293;
  assign T293 = inputReg_2_addr & T294;
  assign T294 = {6'h20/* 32*/{T3}};
  assign T295 = T298 | T296;
  assign T296 = inputReg_1_addr & T297;
  assign T297 = {6'h20/* 32*/{T233}};
  assign T298 = inputReg_0_addr & T299;
  assign T299 = {6'h20/* 32*/{T247}};
  assign T300 = T303 && T301;
  assign T301 = T21 == T302;
  assign T302 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T303 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign mainOff_dram_rep_ready = dramPort_rep_ready;
  assign dramPort_rep_ready = 1'h1/* 1*/;
  assign T304 = ! AllOffloadsReady;
  assign T305 = T350 || T306;
  assign T306 = T346 && T307;
  assign T307 = ! cacheMissPipePort_req_valid;
  assign cacheMissPipePort_req_valid = T308;
  assign T308 = T313 && T309;
  assign T309 = T312 && T310;
  assign T310 = T21 == T311;
  assign T311 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T312 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T313 = T345 && T314;
  assign T314 = ! T315;
  assign T315 = T326 | T316;
  assign T316 = cacheMissPipe_valid_received_2 & T3;
  assign T317 = T323 && T318;
  assign T318 = cacheMissPipe_valid_received_2 || T319;
  assign T319 = cacheMissPipePort_rep_valid && T320;
  assign T320 = cacheMissPipePort_rep_tag == T321;
  assign T321 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign cacheMissPipePort_rep_tag = mainOff_cacheMissPipe_rep_tag;
  assign mainOff_cacheMissPipe_rep_ready = cacheMissPipePort_rep_ready;
  assign cacheMissPipePort_rep_ready = 1'h1/* 1*/;
  assign mainOff_cacheMissPipe_req_tag = cacheMissPipePort_req_tag;
  assign cacheMissPipePort_req_tag = T322;
  assign T322 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign cacheMissPipePort_rep_valid = mainOff_cacheMissPipe_rep_valid;
  assign mainOff_cacheMissPipe_req_valid = cacheMissPipePort_req_valid;
  assign T323 = ! T324;
  assign T324 = T325 == 5'h2/* 2*/;
  assign T325 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T326 = T336 | T327;
  assign T327 = cacheMissPipe_valid_received_1 & T233;
  assign T328 = T333 && T329;
  assign T329 = cacheMissPipe_valid_received_1 || T330;
  assign T330 = cacheMissPipePort_rep_valid && T331;
  assign T331 = cacheMissPipePort_rep_tag == T332;
  assign T332 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T333 = ! T334;
  assign T334 = T335 == 5'h1/* 1*/;
  assign T335 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T336 = cacheMissPipe_valid_received_0 & T247;
  assign T337 = T342 && T338;
  assign T338 = cacheMissPipe_valid_received_0 || T339;
  assign T339 = cacheMissPipePort_rep_valid && T340;
  assign T340 = cacheMissPipePort_rep_tag == T341;
  assign T341 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T346 = ! cacheMissPipePortHadReadyRequest;
  assign T347 = T349 && T348;
  assign T348 = cacheMissPipePortHadReadyRequest || cacheMissPipePort_req_valid;
  assign T349 = ! AllOffloadsReady;
  assign T350 = cacheMissPipePort_req_ready || cacheMissPipe_ready_received;
  assign T351 = T353 && T352;
  assign T352 = cacheMissPipe_ready_received || cacheMissPipePort_req_ready;
  assign cacheMissPipePort_req_ready = mainOff_cacheMissPipe_req_ready;
  assign T353 = ! AllOffloadsReady;
  assign T354 = T396 && T355;
  assign T355 = State_0 == 8'h0/* 0*/;
  assign T356 = T358 || T357;
  assign T357 = T29 && T129;
  assign T358 = T360 || T359;
  assign T359 = T43 && T129;
  assign T360 = T362 || T361;
  assign T361 = T49 && T129;
  assign T362 = T364 || T363;
  assign T363 = T55 && T129;
  assign T364 = T367 || T365;
  assign T365 = T366 && T129;
  assign T366 = T133 && T57;
  assign T367 = T130 || T368;
  assign T368 = T369 && T247;
  assign T369 = T370 && io_out_ready;
  assign T370 = T372 && T371;
  assign T371 = T21 == 8'hff/* 255*/;
  assign T372 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T373 = T357 ? 8'hff/* 255*/ : T374;
  assign T374 = T359 ? T395 : T375;
  assign T375 = T361 ? T394 : T376;
  assign T376 = T363 ? T393 : T377;
  assign T377 = T365 ? T392 : T378;
  assign T378 = T368 ? T381 : T379;
  assign T379 = T130 ? T380 : State_0;
  assign T380 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T381 = T385 | T382;
  assign T382 = EmitReturnState_2 & T383;
  assign T383 = {4'h8/* 8*/{T3}};
  assign T384 = T25 ? 8'h0/* 0*/ : EmitReturnState_2;
  assign T385 = T389 | T386;
  assign T386 = EmitReturnState_1 & T387;
  assign T387 = {4'h8/* 8*/{T233}};
  assign T388 = T40 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T389 = EmitReturnState_0 & T390;
  assign T390 = {4'h8/* 8*/{T247}};
  assign T391 = T357 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T392 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T393 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T394 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T395 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T396 = subStateTh_0 == 1'h0/* 0*/;
  assign T397 = T401 ? 1'h1/* 1*/ : T398;
  assign T398 = T399 ? 1'h0/* 0*/ : subStateTh_0;
  assign T399 = T400 == vThreadEncoder_io_chosen;
  assign T400 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T401 = T403 && T402;
  assign T402 = State_0 != 8'hff/* 255*/;
  assign T403 = T405 && T404;
  assign T404 = State_0 != 8'h0/* 0*/;
  assign T405 = AllOffloadsReady && T406;
  assign T406 = T407 == rThreadEncoder_io_chosen;
  assign T407 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T408 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T409 = T62 ? io_in_bits_rw : inputReg_2_rw;
  assign T410 = T412 | T411;
  assign T411 = inputReg_1_rw & T38;
  assign T412 = inputReg_0_rw & T129;
  assign T413 = ct == T414;
  assign T414 = T421 | T415;
  assign T415 = cachedAddr_2 & T416;
  assign T416 = {6'h20/* 32*/{T26}};
  assign T417 = T62 || T418;
  assign T418 = T55 && T26;
  assign T419 = T418 ? ct : T420;
  assign T420 = T62 ? 32'h0/* 0*/ : cachedAddr_2;
  assign ct = T115 >> 32'h4/* 4*/;
  assign T421 = T427 | T422;
  assign T422 = cachedAddr_1 & T423;
  assign T423 = {6'h20/* 32*/{T38}};
  assign T424 = T122 || T54;
  assign T425 = T54 ? ct : T426;
  assign T426 = T122 ? 32'h0/* 0*/ : cachedAddr_1;
  assign T427 = cachedAddr_0 & T428;
  assign T428 = {6'h20/* 32*/{T129}};
  assign T429 = T130 || T363;
  assign T430 = T363 ? ct : T431;
  assign T431 = T130 ? 32'h0/* 0*/ : cachedAddr_0;
  assign T432 = T434 || T433;
  assign T433 = T366 && T38;
  assign T434 = T122 || T435;
  assign T435 = T369 && T233;
  assign T436 = T40 ? 8'hff/* 255*/ : T437;
  assign T437 = T42 ? T447 : T438;
  assign T438 = T48 ? T446 : T439;
  assign T439 = T54 ? T445 : T440;
  assign T440 = T433 ? T444 : T441;
  assign T441 = T435 ? T381 : T442;
  assign T442 = T122 ? T443 : State_1;
  assign T443 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T444 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T445 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T446 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T447 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T448 = State_0 & T449;
  assign T449 = {4'h8/* 8*/{T129}};
  assign T450 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T451 = T453 || T452;
  assign T452 = T43 && T26;
  assign T453 = T455 || T454;
  assign T454 = T49 && T26;
  assign T455 = T456 || T418;
  assign T456 = T458 || T457;
  assign T457 = T366 && T26;
  assign T458 = T62 || T459;
  assign T459 = T369 && T3;
  assign T460 = T25 ? 8'hff/* 255*/ : T461;
  assign T461 = T452 ? T471 : T462;
  assign T462 = T454 ? T470 : T463;
  assign T463 = T418 ? T469 : T464;
  assign T464 = T457 ? T468 : T465;
  assign T465 = T459 ? T381 : T466;
  assign T466 = T62 ? T467 : State_2;
  assign T467 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T468 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T469 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T470 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T471 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T472 = T475 | T473;
  assign T473 = State_1 & T474;
  assign T474 = {4'h8/* 8*/{T233}};
  assign T475 = State_0 & T476;
  assign T476 = {4'h8/* 8*/{T247}};
  assign T477 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T478 = T510 && T479;
  assign T479 = ! T480;
  assign T480 = T491 | T481;
  assign T481 = dram_valid_received_2 & T3;
  assign T482 = T488 && T483;
  assign T483 = dram_valid_received_2 || T484;
  assign T484 = dramPort_rep_valid && T485;
  assign T485 = dramPort_rep_tag == T486;
  assign T486 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign dramPort_rep_tag = mainOff_dram_rep_tag;
  assign mainOff_dram_req_tag = dramPort_req_tag;
  assign dramPort_req_tag = T487;
  assign T487 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramPort_rep_valid = mainOff_dram_rep_valid;
  assign T488 = ! T489;
  assign T489 = T490 == 5'h2/* 2*/;
  assign T490 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T491 = T501 | T492;
  assign T492 = dram_valid_received_1 & T233;
  assign T493 = T498 && T494;
  assign T494 = dram_valid_received_1 || T495;
  assign T495 = dramPort_rep_valid && T496;
  assign T496 = dramPort_rep_tag == T497;
  assign T497 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T498 = ! T499;
  assign T499 = T500 == 5'h1/* 1*/;
  assign T500 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T501 = dram_valid_received_0 & T247;
  assign T502 = T507 && T503;
  assign T503 = dram_valid_received_0 || T504;
  assign T504 = dramPort_rep_valid && T505;
  assign T505 = dramPort_rep_tag == T506;
  assign T506 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T507 = ! T508;
  assign T508 = T509 == 5'h0/* 0*/;
  assign T509 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T510 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T511 = 5'h2/* 2*/ == T512;
  assign T512 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T513 = ! T514;
  assign T514 = T515 == 5'h2/* 2*/;
  assign T515 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T516 = T517 || dram_valid_received_2;
  assign T517 = dramPort_rep_valid && T518;
  assign T518 = dramPort_rep_tag == T519;
  assign T519 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T520 = T530 || T521;
  assign T521 = ! cacheMissPipePortHadValidRequest_2;
  assign T522 = T527 && T523;
  assign T523 = cacheMissPipePortHadValidRequest_2 || T524;
  assign T524 = T525 && cacheMissPipePort_req_valid;
  assign T525 = 5'h2/* 2*/ == T526;
  assign T526 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T527 = ! T528;
  assign T528 = T529 == 5'h2/* 2*/;
  assign T529 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T530 = T531 || cacheMissPipe_valid_received_2;
  assign T531 = cacheMissPipePort_rep_valid && T532;
  assign T532 = cacheMissPipePort_rep_tag == T533;
  assign T533 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T534 = subStateTh_2 == 1'h1/* 1*/;
  assign T535 = T565 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T536;
  assign T536 = T551 && T537;
  assign T537 = T547 || T538;
  assign T538 = ! dramPortHadValidRequest_1;
  assign T539 = T544 && T540;
  assign T540 = dramPortHadValidRequest_1 || T541;
  assign T541 = T542 && dramPort_req_valid;
  assign T542 = 5'h1/* 1*/ == T543;
  assign T543 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T544 = ! T545;
  assign T545 = T546 == 5'h1/* 1*/;
  assign T546 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T547 = T548 || dram_valid_received_1;
  assign T548 = dramPort_rep_valid && T549;
  assign T549 = dramPort_rep_tag == T550;
  assign T550 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T551 = T561 || T552;
  assign T552 = ! cacheMissPipePortHadValidRequest_1;
  assign T553 = T558 && T554;
  assign T554 = cacheMissPipePortHadValidRequest_1 || T555;
  assign T555 = T556 && cacheMissPipePort_req_valid;
  assign T556 = 5'h1/* 1*/ == T557;
  assign T557 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T558 = ! T559;
  assign T559 = T560 == 5'h1/* 1*/;
  assign T560 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T561 = T562 || cacheMissPipe_valid_received_1;
  assign T562 = cacheMissPipePort_rep_valid && T563;
  assign T563 = cacheMissPipePort_rep_tag == T564;
  assign T564 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T565 = subStateTh_1 == 1'h1/* 1*/;
  assign T566 = T596 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T567;
  assign T567 = T582 && T568;
  assign T568 = T578 || T569;
  assign T569 = ! dramPortHadValidRequest_0;
  assign T570 = T575 && T571;
  assign T571 = dramPortHadValidRequest_0 || T572;
  assign T572 = T573 && dramPort_req_valid;
  assign T573 = 5'h0/* 0*/ == T574;
  assign T574 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T575 = ! T576;
  assign T576 = T577 == 5'h0/* 0*/;
  assign T577 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T578 = T579 || dram_valid_received_0;
  assign T579 = dramPort_rep_valid && T580;
  assign T580 = dramPort_rep_tag == T581;
  assign T581 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T582 = T592 || T583;
  assign T583 = ! cacheMissPipePortHadValidRequest_0;
  assign T584 = T589 && T585;
  assign T585 = cacheMissPipePortHadValidRequest_0 || T586;
  assign T586 = T587 && cacheMissPipePort_req_valid;
  assign T587 = 5'h0/* 0*/ == T588;
  assign T588 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T589 = ! T590;
  assign T590 = T591 == 5'h0/* 0*/;
  assign T591 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T592 = T593 || cacheMissPipe_valid_received_0;
  assign T593 = cacheMissPipePort_rep_valid && T594;
  assign T594 = cacheMissPipePort_rep_tag == T595;
  assign T595 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T596 = subStateTh_0 == 1'h1/* 1*/;
  assign T597 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T598 = T600 && T599;
  assign T599 = State_2 != 8'hff/* 255*/;
  assign T600 = T602 && T601;
  assign T601 = State_2 != 8'h0/* 0*/;
  assign T602 = AllOffloadsReady && T603;
  assign T603 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign T604 = subStateTh_1 == 1'h0/* 0*/;
  assign T605 = subStateTh_0 == 1'h0/* 0*/;
  assign T606 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T607 = T62 ? io_in_tag : inputTag_2;
  assign T608 = T612 | T609;
  assign T609 = inputTag_1 & T610;
  assign T610 = {4'ha/* 10*/{T233}};
  assign T611 = T122 ? io_in_tag : inputTag_1;
  assign T612 = inputTag_0 & T613;
  assign T613 = {4'ha/* 10*/{T247}};
  assign T614 = T130 ? io_in_tag : inputTag_0;
  RREncode_56 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T605 ),
       .io_valid_1( T604 ),
       .io_valid_2( T6 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T606 ));
  RREncode_57 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T566 ),
       .io_valid_1( T535 ),
       .io_valid_2( T10 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T597 ));
  RREncode_58 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T354 ),
       .io_valid_1( T69 ),
       .io_valid_2( T66 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T408 ));

  always @(posedge clk) begin
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T7;
    dramPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T14;
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T24) begin
      State_2 <= T460;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T39) begin
      State_1 <= T436;
    end
    if(T62) begin
      inputReg_2_rw <= T409;
    end
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T72;
    dramPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T88;
    dram_ready_received <= reset ? 1'h0/* 0*/ : T92;
    if(T62) begin
      inputReg_2_size <= T101;
    end
    if(T109) begin
      outputReg_2_data <= T147;
    end
    if(T62) begin
      inputReg_2_addr <= T118;
    end
    if(T122) begin
      inputReg_1_addr <= T126;
    end
    if(T130) begin
      inputReg_0_addr <= T132;
    end
    if(reset) begin
      random_2 <= 32'h1/* 1*/;
    end else if(T158) begin
      random_2 <= T205;
    end
    if(reset) begin
      burst_2 <= 32'h1/* 1*/;
    end else if(T165) begin
      burst_2 <= T173;
    end
    if(reset) begin
      burst_1 <= 32'h1/* 1*/;
    end else if(T180) begin
      burst_1 <= T184;
    end
    if(reset) begin
      burst_0 <= 32'h1/* 1*/;
    end else if(T189) begin
      burst_0 <= T193;
    end
    if(reset) begin
      random_1 <= 32'h1/* 1*/;
    end else if(T212) begin
      random_1 <= T216;
    end
    if(reset) begin
      random_0 <= 32'h1/* 1*/;
    end else if(T221) begin
      random_0 <= T225;
    end
    if(T234) begin
      outputReg_1_data <= T239;
    end
    if(T248) begin
      outputReg_0_data <= T253;
    end
    if(T122) begin
      inputReg_1_size <= T262;
    end
    if(T130) begin
      inputReg_0_size <= T265;
    end
    if(T62) begin
      inputReg_2_data <= T269;
    end
    if(T122) begin
      inputReg_1_data <= T273;
    end
    if(T130) begin
      inputReg_0_data <= T276;
    end
    if(T62) begin
      inputReg_2_cached <= T279;
    end
    if(T122) begin
      inputReg_1_cached <= T282;
    end
    if(T130) begin
      inputReg_0_cached <= T284;
    end
    if(T122) begin
      inputReg_1_rw <= T289;
    end
    if(T130) begin
      inputReg_0_rw <= T291;
    end
    cacheMissPipe_valid_received_2 <= reset ? 1'h0/* 0*/ : T317;
    cacheMissPipe_valid_received_1 <= reset ? 1'h0/* 0*/ : T328;
    cacheMissPipe_valid_received_0 <= reset ? 1'h0/* 0*/ : T337;
    cacheMissPipePortHadReadyRequest <= reset ? 1'h0/* 0*/ : T347;
    cacheMissPipe_ready_received <= reset ? 1'h0/* 0*/ : T351;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T356) begin
      State_0 <= T373;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T25) begin
      EmitReturnState_2 <= T384;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T40) begin
      EmitReturnState_1 <= T388;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T357) begin
      EmitReturnState_0 <= T391;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T397;
    if(reset) begin
      cachedAddr_2 <= 32'h0/* 0*/;
    end else if(T417) begin
      cachedAddr_2 <= T419;
    end
    if(reset) begin
      cachedAddr_1 <= 32'h0/* 0*/;
    end else if(T424) begin
      cachedAddr_1 <= T425;
    end
    if(reset) begin
      cachedAddr_0 <= 32'h0/* 0*/;
    end else if(T429) begin
      cachedAddr_0 <= T430;
    end
    dram_valid_received_2 <= reset ? 1'h0/* 0*/ : T482;
    dram_valid_received_1 <= reset ? 1'h0/* 0*/ : T493;
    dram_valid_received_0 <= reset ? 1'h0/* 0*/ : T502;
    cacheMissPipePortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T522;
    dramPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T539;
    cacheMissPipePortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T553;
    dramPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T570;
    cacheMissPipePortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T584;
    if(T62) begin
      inputTag_2 <= T607;
    end
    if(T122) begin
      inputTag_1 <= T611;
    end
    if(T130) begin
      inputTag_0 <= T614;
    end
  end
endmodule

module gPipe_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_1};
  assign io_out_valid = valids_1;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module gOffloadedComponent_22(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dram_req_ready,
    output mainOff_dram_req_valid,
    output[31:0] mainOff_dram_req_bits_addr,
    output mainOff_dram_req_bits_rw,
    output mainOff_dram_req_bits_cached,
    output[127:0] mainOff_dram_req_bits_data,
    output[3:0] mainOff_dram_req_bits_size,
    output[9:0] mainOff_dram_req_tag,
    output mainOff_dram_rep_ready,
    input  mainOff_dram_rep_valid,
    input [127:0] mainOff_dram_rep_bits_data,
    input [9:0] mainOff_dram_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_dram_req_valid;
  wire[31:0] mainComp_mainOff_dram_req_bits_addr;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[127:0] mainComp_io_out_bits_data;
  wire mainComp_mainOff_dram_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_cacheMissPipe_rep_ready;
  wire[9:0] mainComp_mainOff_cacheMissPipe_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_cacheMissPipe_req_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dram_req_tag;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_dram_req_valid = mainComp_mainOff_dram_req_valid;
  assign mainOff_dram_req_bits_addr = mainComp_mainOff_dram_req_bits_addr;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_bits_data = mainComp_io_out_bits_data;
  assign mainOff_dram_rep_ready = mainComp_mainOff_dram_rep_ready;
  assign mainOff_dram_req_tag = mainComp_mainOff_dram_req_tag;
  cache_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data( mainComp_io_out_bits_data ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_cacheMissPipe_req_ready( offComp_io_in_ready ),
       .mainOff_cacheMissPipe_req_valid( mainComp_mainOff_cacheMissPipe_req_valid ),
       .mainOff_cacheMissPipe_req_bits(  ),
       .mainOff_cacheMissPipe_req_tag( mainComp_mainOff_cacheMissPipe_req_tag ),
       .mainOff_cacheMissPipe_rep_ready( mainComp_mainOff_cacheMissPipe_rep_ready ),
       .mainOff_cacheMissPipe_rep_valid( offComp_io_out_valid ),
       .mainOff_cacheMissPipe_rep_bits(  ),
       .mainOff_cacheMissPipe_rep_tag( offComp_io_out_tag ),
       .mainOff_dram_req_ready( mainOff_dram_req_ready ),
       .mainOff_dram_req_valid( mainComp_mainOff_dram_req_valid ),
       .mainOff_dram_req_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .mainOff_dram_req_bits_rw(  ),
       .mainOff_dram_req_bits_cached(  ),
       .mainOff_dram_req_bits_data(  ),
       .mainOff_dram_req_bits_size(  ),
       .mainOff_dram_req_tag( mainComp_mainOff_dram_req_tag ),
       .mainOff_dram_rep_ready( mainComp_mainOff_dram_rep_ready ),
       .mainOff_dram_rep_valid( mainOff_dram_rep_valid ),
       .mainOff_dram_rep_bits_data(  ),
       .mainOff_dram_rep_tag( mainOff_dram_rep_tag ));
  gPipe_9 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_cacheMissPipe_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_cacheMissPipe_req_tag ),
       .io_out_ready( mainComp_mainOff_cacheMissPipe_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_59(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module RREncode_60(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module RREncode_61(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    input  io_valid_3,
    input  io_valid_4,
    input  io_valid_5,
    input  io_valid_6,
    input  io_valid_7,
    output[3:0] io_chosen,
    input  io_ready);

  wire[3:0] choose;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire T23;
  wire T24;
  reg[2:0] last_grant;
  wire T25;
  wire outValid;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire[2:0] T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[2:0] T54;

  assign io_chosen = choose;
  assign choose = T52 ? T51 : T0;
  assign T0 = T48 ? T47 : T1;
  assign T1 = T44 ? T43 : T2;
  assign T2 = T41 ? T40 : T3;
  assign T3 = T38 ? T37 : T4;
  assign T4 = T35 ? T34 : T5;
  assign T5 = T23 ? T22 : T6;
  assign T6 = io_valid_0 ? T21 : T7;
  assign T7 = io_valid_1 ? T20 : T8;
  assign T8 = io_valid_2 ? T19 : T9;
  assign T9 = io_valid_3 ? T18 : T10;
  assign T10 = io_valid_4 ? T17 : T11;
  assign T11 = io_valid_5 ? T16 : T12;
  assign T12 = io_valid_6 ? T15 : T13;
  assign T13 = io_valid_7 ? T14 : 4'h8/* 8*/;
  assign T14 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T15 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T16 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T17 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T18 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T19 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T20 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T21 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T22 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T23 = io_valid_7 && T24;
  assign T24 = 3'h7/* 7*/ > last_grant;
  assign T25 = outValid && io_ready;
  assign outValid = T26 || io_valid_7;
  assign T26 = T27 || io_valid_6;
  assign T27 = T28 || io_valid_5;
  assign T28 = T29 || io_valid_4;
  assign T29 = T30 || io_valid_3;
  assign T30 = T31 || io_valid_2;
  assign T31 = io_valid_0 || io_valid_1;
  assign T32 = T25 ? choose : T33;
  assign T33 = {1'h0/* 0*/, last_grant};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = io_valid_6 && T36;
  assign T36 = 3'h6/* 6*/ > last_grant;
  assign T37 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = io_valid_5 && T39;
  assign T39 = 3'h5/* 5*/ > last_grant;
  assign T40 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T41 = io_valid_4 && T42;
  assign T42 = 3'h4/* 4*/ > last_grant;
  assign T43 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T44 = io_valid_3 && T45;
  assign T45 = T46 > last_grant;
  assign T46 = {1'h0/* 0*/, 2'h3/* 3*/};
  assign T47 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T48 = io_valid_2 && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 2'h2/* 2*/};
  assign T51 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T52 = io_valid_1 && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {2'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0/* 0*/;
    end else if(T25) begin
      last_grant <= T32;
    end
  end
endmodule

module dram_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank0_req_ready,
    output mainOff_dramBank0_req_valid,
    output[31:0] mainOff_dramBank0_req_bits,
    output[9:0] mainOff_dramBank0_req_tag,
    output mainOff_dramBank0_rep_ready,
    input  mainOff_dramBank0_rep_valid,
    input [31:0] mainOff_dramBank0_rep_bits,
    input [9:0] mainOff_dramBank0_rep_tag,
    input  mainOff_dramBank1_req_ready,
    output mainOff_dramBank1_req_valid,
    output[31:0] mainOff_dramBank1_req_bits,
    output[9:0] mainOff_dramBank1_req_tag,
    output mainOff_dramBank1_rep_ready,
    input  mainOff_dramBank1_rep_valid,
    input [31:0] mainOff_dramBank1_rep_bits,
    input [9:0] mainOff_dramBank1_rep_tag,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire T0;
  wire[3:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_7;
  wire T3;
  wire T4;
  wire T5;
  wire[7:0] T6;
  wire[22:0] T7;
  wire[3:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_7;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] dramBank7PortHadValidRequest_7;
  wire T12;
  wire T13;
  wire T14;
  wire dramBank7Port_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire[7:0] T23;
  wire[22:0] T24;
  wire[3:0] rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_7;
  wire T26;
  wire T27;
  wire T28;
  wire[3:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[3:0] T36;
  wire AllOffloadsReady;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg[0:0] dramBank7PortHadReadyRequest;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  reg[0:0] dramBank7_ready_received;
  wire T46;
  wire T47;
  wire dramBank7Port_req_ready;
  wire dramBank7Port_rep_ready;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire dramBank6Port_req_valid;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  reg[0:0] dramBank6_valid_received_7;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[9:0] T66;
  wire[9:0] dramBank6Port_rep_tag;
  wire dramBank6Port_rep_ready;
  wire[9:0] dramBank6Port_req_tag;
  wire[9:0] T67;
  wire dramBank6Port_rep_valid;
  wire T68;
  wire T69;
  wire[4:0] T70;
  wire T71;
  wire T72;
  wire T73;
  reg[0:0] dramBank6_valid_received_6;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[9:0] T78;
  wire T79;
  wire T80;
  wire[4:0] T81;
  wire T82;
  wire T83;
  wire T84;
  reg[0:0] dramBank6_valid_received_5;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire[9:0] T89;
  wire T90;
  wire T91;
  wire[4:0] T92;
  wire T93;
  wire T94;
  wire T95;
  reg[0:0] dramBank6_valid_received_4;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[9:0] T100;
  wire T101;
  wire T102;
  wire[4:0] T103;
  wire T104;
  wire T105;
  wire T106;
  reg[0:0] dramBank6_valid_received_3;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[9:0] T111;
  wire T112;
  wire T113;
  wire[4:0] T114;
  wire T115;
  wire T116;
  wire T117;
  reg[0:0] dramBank6_valid_received_2;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[9:0] T122;
  wire T123;
  wire T124;
  wire[4:0] T125;
  wire T126;
  wire T127;
  wire T128;
  reg[0:0] dramBank6_valid_received_1;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire[9:0] T133;
  wire T134;
  wire T135;
  wire[4:0] T136;
  wire T137;
  wire T138;
  reg[0:0] dramBank6_valid_received_0;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire[9:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  reg[0:0] dramBank6PortHadReadyRequest;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] dramBank6_ready_received;
  wire T153;
  wire T154;
  wire dramBank6Port_req_ready;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire dramBank5Port_req_valid;
  wire T160;
  wire T161;
  wire T162;
  wire[7:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  reg[0:0] dramBank5_valid_received_7;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[9:0] T173;
  wire[9:0] dramBank5Port_rep_tag;
  wire dramBank5Port_rep_ready;
  wire[9:0] dramBank5Port_req_tag;
  wire[9:0] T174;
  wire dramBank5Port_rep_valid;
  wire T175;
  wire T176;
  wire[4:0] T177;
  wire T178;
  wire T179;
  reg[0:0] dramBank5_valid_received_6;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[9:0] T184;
  wire T185;
  wire T186;
  wire[4:0] T187;
  wire T188;
  wire T189;
  reg[0:0] dramBank5_valid_received_5;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire[9:0] T194;
  wire T195;
  wire T196;
  wire[4:0] T197;
  wire T198;
  wire T199;
  reg[0:0] dramBank5_valid_received_4;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[9:0] T204;
  wire T205;
  wire T206;
  wire[4:0] T207;
  wire T208;
  wire T209;
  reg[0:0] dramBank5_valid_received_3;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[9:0] T214;
  wire T215;
  wire T216;
  wire[4:0] T217;
  wire T218;
  wire T219;
  reg[0:0] dramBank5_valid_received_2;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[9:0] T224;
  wire T225;
  wire T226;
  wire[4:0] T227;
  wire T228;
  wire T229;
  reg[0:0] dramBank5_valid_received_1;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire[9:0] T234;
  wire T235;
  wire T236;
  wire[4:0] T237;
  wire T238;
  reg[0:0] dramBank5_valid_received_0;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire[9:0] T243;
  wire T244;
  wire T245;
  wire[4:0] T246;
  wire T247;
  wire T248;
  reg[0:0] dramBank5PortHadReadyRequest;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] dramBank5_ready_received;
  wire T253;
  wire T254;
  wire dramBank5Port_req_ready;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire dramBank4Port_req_valid;
  wire T260;
  wire T261;
  wire T262;
  wire[7:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  reg[0:0] dramBank4_valid_received_7;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[9:0] T273;
  wire[9:0] dramBank4Port_rep_tag;
  wire dramBank4Port_rep_ready;
  wire[9:0] dramBank4Port_req_tag;
  wire[9:0] T274;
  wire dramBank4Port_rep_valid;
  wire T275;
  wire T276;
  wire[4:0] T277;
  wire T278;
  wire T279;
  reg[0:0] dramBank4_valid_received_6;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[9:0] T284;
  wire T285;
  wire T286;
  wire[4:0] T287;
  wire T288;
  wire T289;
  reg[0:0] dramBank4_valid_received_5;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[9:0] T294;
  wire T295;
  wire T296;
  wire[4:0] T297;
  wire T298;
  wire T299;
  reg[0:0] dramBank4_valid_received_4;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[9:0] T304;
  wire T305;
  wire T306;
  wire[4:0] T307;
  wire T308;
  wire T309;
  reg[0:0] dramBank4_valid_received_3;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire[9:0] T314;
  wire T315;
  wire T316;
  wire[4:0] T317;
  wire T318;
  wire T319;
  reg[0:0] dramBank4_valid_received_2;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[9:0] T324;
  wire T325;
  wire T326;
  wire[4:0] T327;
  wire T328;
  wire T329;
  reg[0:0] dramBank4_valid_received_1;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire T335;
  wire T336;
  wire[4:0] T337;
  wire T338;
  reg[0:0] dramBank4_valid_received_0;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire[9:0] T343;
  wire T344;
  wire T345;
  wire[4:0] T346;
  wire T347;
  wire T348;
  reg[0:0] dramBank4PortHadReadyRequest;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  reg[0:0] dramBank4_ready_received;
  wire T353;
  wire T354;
  wire dramBank4Port_req_ready;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire dramBank3Port_req_valid;
  wire T360;
  wire T361;
  wire T362;
  wire[7:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  reg[0:0] dramBank3_valid_received_7;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire[9:0] T373;
  wire[9:0] dramBank3Port_rep_tag;
  wire dramBank3Port_rep_ready;
  wire[9:0] dramBank3Port_req_tag;
  wire[9:0] T374;
  wire dramBank3Port_rep_valid;
  wire T375;
  wire T376;
  wire[4:0] T377;
  wire T378;
  wire T379;
  reg[0:0] dramBank3_valid_received_6;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire[9:0] T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire T388;
  wire T389;
  reg[0:0] dramBank3_valid_received_5;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[9:0] T394;
  wire T395;
  wire T396;
  wire[4:0] T397;
  wire T398;
  wire T399;
  reg[0:0] dramBank3_valid_received_4;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[9:0] T404;
  wire T405;
  wire T406;
  wire[4:0] T407;
  wire T408;
  wire T409;
  reg[0:0] dramBank3_valid_received_3;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire[9:0] T414;
  wire T415;
  wire T416;
  wire[4:0] T417;
  wire T418;
  wire T419;
  reg[0:0] dramBank3_valid_received_2;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[9:0] T424;
  wire T425;
  wire T426;
  wire[4:0] T427;
  wire T428;
  wire T429;
  reg[0:0] dramBank3_valid_received_1;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire[9:0] T434;
  wire T435;
  wire T436;
  wire[4:0] T437;
  wire T438;
  reg[0:0] dramBank3_valid_received_0;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire[9:0] T443;
  wire T444;
  wire T445;
  wire[4:0] T446;
  wire T447;
  wire T448;
  reg[0:0] dramBank3PortHadReadyRequest;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] dramBank3_ready_received;
  wire T453;
  wire T454;
  wire dramBank3Port_req_ready;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire dramBank2Port_req_valid;
  wire T460;
  wire T461;
  wire T462;
  wire[7:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] dramBank2_valid_received_7;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire[9:0] T473;
  wire[9:0] dramBank2Port_rep_tag;
  wire dramBank2Port_rep_ready;
  wire[9:0] dramBank2Port_req_tag;
  wire[9:0] T474;
  wire dramBank2Port_rep_valid;
  wire T475;
  wire T476;
  wire[4:0] T477;
  wire T478;
  wire T479;
  reg[0:0] dramBank2_valid_received_6;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[9:0] T484;
  wire T485;
  wire T486;
  wire[4:0] T487;
  wire T488;
  wire T489;
  reg[0:0] dramBank2_valid_received_5;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[9:0] T494;
  wire T495;
  wire T496;
  wire[4:0] T497;
  wire T498;
  wire T499;
  reg[0:0] dramBank2_valid_received_4;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[9:0] T504;
  wire T505;
  wire T506;
  wire[4:0] T507;
  wire T508;
  wire T509;
  reg[0:0] dramBank2_valid_received_3;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire[9:0] T514;
  wire T515;
  wire T516;
  wire[4:0] T517;
  wire T518;
  wire T519;
  reg[0:0] dramBank2_valid_received_2;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[9:0] T524;
  wire T525;
  wire T526;
  wire[4:0] T527;
  wire T528;
  wire T529;
  reg[0:0] dramBank2_valid_received_1;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[9:0] T534;
  wire T535;
  wire T536;
  wire[4:0] T537;
  wire T538;
  reg[0:0] dramBank2_valid_received_0;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire[9:0] T543;
  wire T544;
  wire T545;
  wire[4:0] T546;
  wire T547;
  wire T548;
  reg[0:0] dramBank2PortHadReadyRequest;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  reg[0:0] dramBank2_ready_received;
  wire T553;
  wire T554;
  wire dramBank2Port_req_ready;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire dramBank1Port_req_valid;
  wire T560;
  wire T561;
  wire T562;
  wire[7:0] T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  reg[0:0] dramBank1_valid_received_7;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire[9:0] T573;
  wire[9:0] dramBank1Port_rep_tag;
  wire dramBank1Port_rep_ready;
  wire[9:0] dramBank1Port_req_tag;
  wire[9:0] T574;
  wire dramBank1Port_rep_valid;
  wire T575;
  wire T576;
  wire[4:0] T577;
  wire T578;
  wire T579;
  reg[0:0] dramBank1_valid_received_6;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire[9:0] T584;
  wire T585;
  wire T586;
  wire[4:0] T587;
  wire T588;
  wire T589;
  reg[0:0] dramBank1_valid_received_5;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire[9:0] T594;
  wire T595;
  wire T596;
  wire[4:0] T597;
  wire T598;
  wire T599;
  reg[0:0] dramBank1_valid_received_4;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[9:0] T604;
  wire T605;
  wire T606;
  wire[4:0] T607;
  wire T608;
  wire T609;
  reg[0:0] dramBank1_valid_received_3;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[9:0] T614;
  wire T615;
  wire T616;
  wire[4:0] T617;
  wire T618;
  wire T619;
  reg[0:0] dramBank1_valid_received_2;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[9:0] T624;
  wire T625;
  wire T626;
  wire[4:0] T627;
  wire T628;
  wire T629;
  reg[0:0] dramBank1_valid_received_1;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire[9:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  reg[0:0] dramBank1_valid_received_0;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire[9:0] T643;
  wire T644;
  wire T645;
  wire[4:0] T646;
  wire T647;
  wire T648;
  reg[0:0] dramBank1PortHadReadyRequest;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  reg[0:0] dramBank1_ready_received;
  wire T653;
  wire T654;
  wire dramBank1Port_req_ready;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire dramBank0Port_req_valid;
  wire T659;
  wire T660;
  wire T661;
  wire[7:0] T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  reg[0:0] dramBank0_valid_received_7;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire[9:0] T672;
  wire[9:0] dramBank0Port_rep_tag;
  wire dramBank0Port_rep_ready;
  wire[9:0] dramBank0Port_req_tag;
  wire[9:0] T673;
  wire dramBank0Port_rep_valid;
  wire T674;
  wire T675;
  wire[4:0] T676;
  wire T677;
  wire T678;
  reg[0:0] dramBank0_valid_received_6;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire[9:0] T683;
  wire T684;
  wire T685;
  wire[4:0] T686;
  wire T687;
  wire T688;
  reg[0:0] dramBank0_valid_received_5;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire[9:0] T693;
  wire T694;
  wire T695;
  wire[4:0] T696;
  wire T697;
  wire T698;
  reg[0:0] dramBank0_valid_received_4;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire[9:0] T703;
  wire T704;
  wire T705;
  wire[4:0] T706;
  wire T707;
  wire T708;
  reg[0:0] dramBank0_valid_received_3;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[9:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  reg[0:0] dramBank0_valid_received_2;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire[9:0] T723;
  wire T724;
  wire T725;
  wire[4:0] T726;
  wire T727;
  wire T728;
  reg[0:0] dramBank0_valid_received_1;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire[9:0] T733;
  wire T734;
  wire T735;
  wire[4:0] T736;
  wire T737;
  reg[0:0] dramBank0_valid_received_0;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[9:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  reg[0:0] dramBank0PortHadReadyRequest;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  reg[0:0] dramBank0_ready_received;
  wire T752;
  wire T753;
  wire dramBank0Port_req_ready;
  wire T754;
  wire T755;
  reg[0:0] subStateTh_6;
  wire T756;
  wire T757;
  wire T758;
  wire[3:0] T759;
  wire T760;
  wire T761;
  reg[7:0] State_6;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[7:0] T767;
  wire[7:0] T768;
  wire[7:0] T769;
  wire[7:0] T770;
  wire[7:0] T771;
  wire[7:0] T772;
  wire[7:0] T773;
  wire[7:0] T774;
  wire[7:0] T775;
  wire[7:0] T776;
  wire T777;
  reg[7:0] State_5;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[7:0] T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[7:0] T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[7:0] T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire[7:0] T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire[7:0] T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[7:0] T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[7:0] T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire[7:0] T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire[47:0] T833;
  wire[47:0] b;
  wire[47:0] T834;
  wire[31:0] T835;
  wire[31:0] T836;
  wire[31:0] T837;
  wire[31:0] T838;
  reg[31:0] inputReg_7_addr;
  wire T839;
  wire T840;
  wire[7:0] T841;
  wire[22:0] T842;
  wire T843;
  wire T844;
  wire[31:0] T845;
  wire[31:0] T846;
  wire[31:0] T847;
  wire[31:0] T848;
  reg[31:0] inputReg_6_addr;
  wire T849;
  wire T850;
  wire[31:0] T851;
  wire[31:0] T852;
  wire[31:0] T853;
  wire[31:0] T854;
  reg[31:0] inputReg_5_addr;
  wire T855;
  wire T856;
  wire[31:0] T857;
  wire[31:0] T858;
  wire[31:0] T859;
  wire[31:0] T860;
  wire T861;
  reg[31:0] inputReg_4_addr;
  wire T862;
  wire T863;
  wire[31:0] T864;
  wire[31:0] T865;
  wire[31:0] T866;
  wire[31:0] T867;
  wire T868;
  reg[31:0] inputReg_3_addr;
  wire T869;
  wire T870;
  wire[31:0] T871;
  wire[31:0] T872;
  wire[31:0] T873;
  wire[31:0] T874;
  wire T875;
  reg[31:0] inputReg_2_addr;
  wire T876;
  wire T877;
  wire[31:0] T878;
  wire[31:0] T879;
  wire[31:0] T880;
  wire[31:0] T881;
  wire T882;
  reg[31:0] inputReg_1_addr;
  wire T883;
  wire T884;
  wire[31:0] T885;
  wire[31:0] T886;
  wire[31:0] T887;
  wire T888;
  reg[31:0] inputReg_0_addr;
  wire T889;
  wire T890;
  wire[31:0] T891;
  wire T892;
  wire T893;
  wire T894;
  wire[47:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[47:0] T899;
  wire T900;
  wire T901;
  wire T902;
  wire[47:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[47:0] T907;
  wire T908;
  wire T909;
  wire T910;
  wire[47:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[47:0] T915;
  wire T916;
  wire T917;
  wire T918;
  wire[47:0] T919;
  wire T920;
  wire T921;
  wire[7:0] T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire T928;
  wire[59:0] r;
  wire[59:0] T929;
  wire[31:0] T930;
  wire[59:0] T931;
  wire[31:0] T932;
  wire[31:0] T933;
  wire[31:0] T934;
  reg[31:0] rb7RowAddr_7;
  wire T935;
  wire T936;
  wire[59:0] T937;
  wire[59:0] T938;
  wire[31:0] T939;
  wire[31:0] T940;
  wire[31:0] T941;
  wire[31:0] T942;
  reg[31:0] rb7RowAddr_6;
  wire T943;
  wire T944;
  wire[59:0] T945;
  wire[59:0] T946;
  wire[31:0] T947;
  wire[31:0] T948;
  wire[31:0] T949;
  wire[31:0] T950;
  reg[31:0] rb7RowAddr_5;
  wire T951;
  wire[59:0] T952;
  wire[59:0] T953;
  wire[31:0] T954;
  wire[31:0] T955;
  wire[31:0] T956;
  wire[31:0] T957;
  reg[31:0] rb7RowAddr_4;
  wire T958;
  wire T959;
  wire[59:0] T960;
  wire[59:0] T961;
  wire[31:0] T962;
  wire[31:0] T963;
  wire[31:0] T964;
  wire[31:0] T965;
  reg[31:0] rb7RowAddr_3;
  wire T966;
  wire T967;
  wire[59:0] T968;
  wire[59:0] T969;
  wire[31:0] T970;
  wire[31:0] T971;
  wire[31:0] T972;
  wire[31:0] T973;
  reg[31:0] rb7RowAddr_2;
  wire T974;
  wire T975;
  wire[59:0] T976;
  wire[59:0] T977;
  wire[31:0] T978;
  wire[31:0] T979;
  wire[31:0] T980;
  wire[31:0] T981;
  reg[31:0] rb7RowAddr_1;
  wire T982;
  wire T983;
  wire[59:0] T984;
  wire[59:0] T985;
  wire[31:0] T986;
  wire[31:0] T987;
  wire[31:0] T988;
  reg[31:0] rb7RowAddr_0;
  wire T989;
  wire T990;
  wire[59:0] T991;
  wire[59:0] T992;
  wire[31:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[59:0] T1003;
  wire[31:0] T1004;
  wire[31:0] T1005;
  wire[31:0] T1006;
  reg[31:0] rb6RowAddr_7;
  wire T1007;
  wire T1008;
  wire[59:0] T1009;
  wire[59:0] T1010;
  wire[31:0] T1011;
  wire[31:0] T1012;
  wire[31:0] T1013;
  wire[31:0] T1014;
  reg[31:0] rb6RowAddr_6;
  wire T1015;
  wire T1016;
  wire[59:0] T1017;
  wire[59:0] T1018;
  wire[31:0] T1019;
  wire[31:0] T1020;
  wire[31:0] T1021;
  wire[31:0] T1022;
  reg[31:0] rb6RowAddr_5;
  wire T1023;
  wire[59:0] T1024;
  wire[59:0] T1025;
  wire[31:0] T1026;
  wire[31:0] T1027;
  wire[31:0] T1028;
  wire[31:0] T1029;
  reg[31:0] rb6RowAddr_4;
  wire T1030;
  wire T1031;
  wire[59:0] T1032;
  wire[59:0] T1033;
  wire[31:0] T1034;
  wire[31:0] T1035;
  wire[31:0] T1036;
  wire[31:0] T1037;
  reg[31:0] rb6RowAddr_3;
  wire T1038;
  wire T1039;
  wire[59:0] T1040;
  wire[59:0] T1041;
  wire[31:0] T1042;
  wire[31:0] T1043;
  wire[31:0] T1044;
  wire[31:0] T1045;
  reg[31:0] rb6RowAddr_2;
  wire T1046;
  wire T1047;
  wire[59:0] T1048;
  wire[59:0] T1049;
  wire[31:0] T1050;
  wire[31:0] T1051;
  wire[31:0] T1052;
  wire[31:0] T1053;
  reg[31:0] rb6RowAddr_1;
  wire T1054;
  wire T1055;
  wire[59:0] T1056;
  wire[59:0] T1057;
  wire[31:0] T1058;
  wire[31:0] T1059;
  wire[31:0] T1060;
  reg[31:0] rb6RowAddr_0;
  wire T1061;
  wire T1062;
  wire[59:0] T1063;
  wire[59:0] T1064;
  wire[31:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire[59:0] T1075;
  wire[31:0] T1076;
  wire[31:0] T1077;
  wire[31:0] T1078;
  reg[31:0] rb5RowAddr_7;
  wire T1079;
  wire T1080;
  wire[59:0] T1081;
  wire[59:0] T1082;
  wire[31:0] T1083;
  wire[31:0] T1084;
  wire[31:0] T1085;
  wire[31:0] T1086;
  reg[31:0] rb5RowAddr_6;
  wire T1087;
  wire T1088;
  wire[59:0] T1089;
  wire[59:0] T1090;
  wire[31:0] T1091;
  wire[31:0] T1092;
  wire[31:0] T1093;
  wire[31:0] T1094;
  reg[31:0] rb5RowAddr_5;
  wire T1095;
  wire[59:0] T1096;
  wire[59:0] T1097;
  wire[31:0] T1098;
  wire[31:0] T1099;
  wire[31:0] T1100;
  wire[31:0] T1101;
  reg[31:0] rb5RowAddr_4;
  wire T1102;
  wire T1103;
  wire[59:0] T1104;
  wire[59:0] T1105;
  wire[31:0] T1106;
  wire[31:0] T1107;
  wire[31:0] T1108;
  wire[31:0] T1109;
  reg[31:0] rb5RowAddr_3;
  wire T1110;
  wire T1111;
  wire[59:0] T1112;
  wire[59:0] T1113;
  wire[31:0] T1114;
  wire[31:0] T1115;
  wire[31:0] T1116;
  wire[31:0] T1117;
  reg[31:0] rb5RowAddr_2;
  wire T1118;
  wire T1119;
  wire[59:0] T1120;
  wire[59:0] T1121;
  wire[31:0] T1122;
  wire[31:0] T1123;
  wire[31:0] T1124;
  wire[31:0] T1125;
  reg[31:0] rb5RowAddr_1;
  wire T1126;
  wire T1127;
  wire[59:0] T1128;
  wire[59:0] T1129;
  wire[31:0] T1130;
  wire[31:0] T1131;
  wire[31:0] T1132;
  reg[31:0] rb5RowAddr_0;
  wire T1133;
  wire T1134;
  wire[59:0] T1135;
  wire[59:0] T1136;
  wire[31:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire[59:0] T1147;
  wire[31:0] T1148;
  wire[31:0] T1149;
  wire[31:0] T1150;
  reg[31:0] rb4RowAddr_7;
  wire T1151;
  wire T1152;
  wire[59:0] T1153;
  wire[59:0] T1154;
  wire[31:0] T1155;
  wire[31:0] T1156;
  wire[31:0] T1157;
  wire[31:0] T1158;
  reg[31:0] rb4RowAddr_6;
  wire T1159;
  wire T1160;
  wire[59:0] T1161;
  wire[59:0] T1162;
  wire[31:0] T1163;
  wire[31:0] T1164;
  wire[31:0] T1165;
  wire[31:0] T1166;
  reg[31:0] rb4RowAddr_5;
  wire T1167;
  wire[59:0] T1168;
  wire[59:0] T1169;
  wire[31:0] T1170;
  wire[31:0] T1171;
  wire[31:0] T1172;
  wire[31:0] T1173;
  reg[31:0] rb4RowAddr_4;
  wire T1174;
  wire T1175;
  wire[59:0] T1176;
  wire[59:0] T1177;
  wire[31:0] T1178;
  wire[31:0] T1179;
  wire[31:0] T1180;
  wire[31:0] T1181;
  reg[31:0] rb4RowAddr_3;
  wire T1182;
  wire T1183;
  wire[59:0] T1184;
  wire[59:0] T1185;
  wire[31:0] T1186;
  wire[31:0] T1187;
  wire[31:0] T1188;
  wire[31:0] T1189;
  reg[31:0] rb4RowAddr_2;
  wire T1190;
  wire T1191;
  wire[59:0] T1192;
  wire[59:0] T1193;
  wire[31:0] T1194;
  wire[31:0] T1195;
  wire[31:0] T1196;
  wire[31:0] T1197;
  reg[31:0] rb4RowAddr_1;
  wire T1198;
  wire T1199;
  wire[59:0] T1200;
  wire[59:0] T1201;
  wire[31:0] T1202;
  wire[31:0] T1203;
  wire[31:0] T1204;
  reg[31:0] rb4RowAddr_0;
  wire T1205;
  wire T1206;
  wire[59:0] T1207;
  wire[59:0] T1208;
  wire[31:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire[59:0] T1219;
  wire[31:0] T1220;
  wire[31:0] T1221;
  wire[31:0] T1222;
  reg[31:0] rb3RowAddr_7;
  wire T1223;
  wire T1224;
  wire[59:0] T1225;
  wire[59:0] T1226;
  wire[31:0] T1227;
  wire[31:0] T1228;
  wire[31:0] T1229;
  wire[31:0] T1230;
  reg[31:0] rb3RowAddr_6;
  wire T1231;
  wire T1232;
  wire[59:0] T1233;
  wire[59:0] T1234;
  wire[31:0] T1235;
  wire[31:0] T1236;
  wire[31:0] T1237;
  wire[31:0] T1238;
  reg[31:0] rb3RowAddr_5;
  wire T1239;
  wire[59:0] T1240;
  wire[59:0] T1241;
  wire[31:0] T1242;
  wire[31:0] T1243;
  wire[31:0] T1244;
  wire[31:0] T1245;
  reg[31:0] rb3RowAddr_4;
  wire T1246;
  wire T1247;
  wire[59:0] T1248;
  wire[59:0] T1249;
  wire[31:0] T1250;
  wire[31:0] T1251;
  wire[31:0] T1252;
  wire[31:0] T1253;
  reg[31:0] rb3RowAddr_3;
  wire T1254;
  wire T1255;
  wire[59:0] T1256;
  wire[59:0] T1257;
  wire[31:0] T1258;
  wire[31:0] T1259;
  wire[31:0] T1260;
  wire[31:0] T1261;
  reg[31:0] rb3RowAddr_2;
  wire T1262;
  wire T1263;
  wire[59:0] T1264;
  wire[59:0] T1265;
  wire[31:0] T1266;
  wire[31:0] T1267;
  wire[31:0] T1268;
  wire[31:0] T1269;
  reg[31:0] rb3RowAddr_1;
  wire T1270;
  wire T1271;
  wire[59:0] T1272;
  wire[59:0] T1273;
  wire[31:0] T1274;
  wire[31:0] T1275;
  wire[31:0] T1276;
  reg[31:0] rb3RowAddr_0;
  wire T1277;
  wire T1278;
  wire[59:0] T1279;
  wire[59:0] T1280;
  wire[31:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire[59:0] T1291;
  wire[31:0] T1292;
  wire[31:0] T1293;
  wire[31:0] T1294;
  reg[31:0] rb2RowAddr_7;
  wire T1295;
  wire T1296;
  wire[59:0] T1297;
  wire[59:0] T1298;
  wire[31:0] T1299;
  wire[31:0] T1300;
  wire[31:0] T1301;
  wire[31:0] T1302;
  reg[31:0] rb2RowAddr_6;
  wire T1303;
  wire T1304;
  wire[59:0] T1305;
  wire[59:0] T1306;
  wire[31:0] T1307;
  wire[31:0] T1308;
  wire[31:0] T1309;
  wire[31:0] T1310;
  reg[31:0] rb2RowAddr_5;
  wire T1311;
  wire[59:0] T1312;
  wire[59:0] T1313;
  wire[31:0] T1314;
  wire[31:0] T1315;
  wire[31:0] T1316;
  wire[31:0] T1317;
  reg[31:0] rb2RowAddr_4;
  wire T1318;
  wire T1319;
  wire[59:0] T1320;
  wire[59:0] T1321;
  wire[31:0] T1322;
  wire[31:0] T1323;
  wire[31:0] T1324;
  wire[31:0] T1325;
  reg[31:0] rb2RowAddr_3;
  wire T1326;
  wire T1327;
  wire[59:0] T1328;
  wire[59:0] T1329;
  wire[31:0] T1330;
  wire[31:0] T1331;
  wire[31:0] T1332;
  wire[31:0] T1333;
  reg[31:0] rb2RowAddr_2;
  wire T1334;
  wire T1335;
  wire[59:0] T1336;
  wire[59:0] T1337;
  wire[31:0] T1338;
  wire[31:0] T1339;
  wire[31:0] T1340;
  wire[31:0] T1341;
  reg[31:0] rb2RowAddr_1;
  wire T1342;
  wire T1343;
  wire[59:0] T1344;
  wire[59:0] T1345;
  wire[31:0] T1346;
  wire[31:0] T1347;
  wire[31:0] T1348;
  reg[31:0] rb2RowAddr_0;
  wire T1349;
  wire T1350;
  wire[59:0] T1351;
  wire[59:0] T1352;
  wire[31:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire[59:0] T1363;
  wire[31:0] T1364;
  wire[31:0] T1365;
  wire[31:0] T1366;
  reg[31:0] rb1RowAddr_7;
  wire T1367;
  wire T1368;
  wire[59:0] T1369;
  wire[59:0] T1370;
  wire[31:0] T1371;
  wire[31:0] T1372;
  wire[31:0] T1373;
  wire[31:0] T1374;
  reg[31:0] rb1RowAddr_6;
  wire T1375;
  wire T1376;
  wire[59:0] T1377;
  wire[59:0] T1378;
  wire[31:0] T1379;
  wire[31:0] T1380;
  wire[31:0] T1381;
  wire[31:0] T1382;
  reg[31:0] rb1RowAddr_5;
  wire T1383;
  wire[59:0] T1384;
  wire[59:0] T1385;
  wire[31:0] T1386;
  wire[31:0] T1387;
  wire[31:0] T1388;
  wire[31:0] T1389;
  reg[31:0] rb1RowAddr_4;
  wire T1390;
  wire T1391;
  wire[59:0] T1392;
  wire[59:0] T1393;
  wire[31:0] T1394;
  wire[31:0] T1395;
  wire[31:0] T1396;
  wire[31:0] T1397;
  reg[31:0] rb1RowAddr_3;
  wire T1398;
  wire T1399;
  wire[59:0] T1400;
  wire[59:0] T1401;
  wire[31:0] T1402;
  wire[31:0] T1403;
  wire[31:0] T1404;
  wire[31:0] T1405;
  reg[31:0] rb1RowAddr_2;
  wire T1406;
  wire T1407;
  wire[59:0] T1408;
  wire[59:0] T1409;
  wire[31:0] T1410;
  wire[31:0] T1411;
  wire[31:0] T1412;
  wire[31:0] T1413;
  reg[31:0] rb1RowAddr_1;
  wire T1414;
  wire T1415;
  wire[59:0] T1416;
  wire[59:0] T1417;
  wire[31:0] T1418;
  wire[31:0] T1419;
  wire[31:0] T1420;
  reg[31:0] rb1RowAddr_0;
  wire T1421;
  wire T1422;
  wire[59:0] T1423;
  wire[59:0] T1424;
  wire[31:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire[59:0] T1435;
  wire[31:0] T1436;
  wire[31:0] T1437;
  wire[31:0] T1438;
  reg[31:0] rb0RowAddr_7;
  wire T1439;
  wire T1440;
  wire[59:0] T1441;
  wire[59:0] T1442;
  wire[31:0] T1443;
  wire[31:0] T1444;
  wire[31:0] T1445;
  wire[31:0] T1446;
  reg[31:0] rb0RowAddr_6;
  wire T1447;
  wire T1448;
  wire[59:0] T1449;
  wire[59:0] T1450;
  wire[31:0] T1451;
  wire[31:0] T1452;
  wire[31:0] T1453;
  wire[31:0] T1454;
  reg[31:0] rb0RowAddr_5;
  wire T1455;
  wire[59:0] T1456;
  wire[59:0] T1457;
  wire[31:0] T1458;
  wire[31:0] T1459;
  wire[31:0] T1460;
  wire[31:0] T1461;
  reg[31:0] rb0RowAddr_4;
  wire T1462;
  wire T1463;
  wire[59:0] T1464;
  wire[59:0] T1465;
  wire[31:0] T1466;
  wire[31:0] T1467;
  wire[31:0] T1468;
  wire[31:0] T1469;
  reg[31:0] rb0RowAddr_3;
  wire T1470;
  wire T1471;
  wire[59:0] T1472;
  wire[59:0] T1473;
  wire[31:0] T1474;
  wire[31:0] T1475;
  wire[31:0] T1476;
  wire[31:0] T1477;
  reg[31:0] rb0RowAddr_2;
  wire T1478;
  wire T1479;
  wire[59:0] T1480;
  wire[59:0] T1481;
  wire[31:0] T1482;
  wire[31:0] T1483;
  wire[31:0] T1484;
  wire[31:0] T1485;
  reg[31:0] rb0RowAddr_1;
  wire T1486;
  wire T1487;
  wire[59:0] T1488;
  wire[59:0] T1489;
  wire[31:0] T1490;
  wire[31:0] T1491;
  wire[31:0] T1492;
  reg[31:0] rb0RowAddr_0;
  wire T1493;
  wire T1494;
  wire[59:0] T1495;
  wire[59:0] T1496;
  wire[31:0] T1497;
  wire T1498;
  wire T1499;
  wire T1500;
  wire T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire[7:0] T1508;
  wire[7:0] T1509;
  wire[7:0] T1510;
  wire[7:0] T1511;
  wire[7:0] T1512;
  wire[7:0] T1513;
  wire[7:0] T1514;
  wire[7:0] T1515;
  wire[7:0] T1516;
  wire[7:0] T1517;
  wire[7:0] T1518;
  wire[7:0] T1519;
  wire[7:0] T1520;
  wire[7:0] T1521;
  wire[7:0] T1522;
  wire[7:0] T1523;
  wire[7:0] T1524;
  wire[7:0] T1525;
  wire[7:0] T1526;
  wire[7:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[7:0] T1530;
  wire[7:0] T1531;
  reg[7:0] EmitReturnState_7;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire T1540;
  wire T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  wire T1546;
  wire T1547;
  wire[7:0] T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire T1556;
  wire[7:0] T1557;
  wire[7:0] T1558;
  wire[7:0] T1559;
  reg[7:0] EmitReturnState_6;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire T1564;
  wire T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire[7:0] T1576;
  wire T1577;
  wire T1578;
  wire T1579;
  wire T1580;
  wire T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[7:0] T1585;
  wire[7:0] T1586;
  wire[7:0] T1587;
  reg[7:0] EmitReturnState_5;
  wire T1588;
  wire T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire[7:0] T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire T1604;
  wire[7:0] T1605;
  wire[7:0] T1606;
  wire[7:0] T1607;
  reg[7:0] EmitReturnState_4;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire T1620;
  wire T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[7:0] T1625;
  wire T1626;
  wire T1627;
  wire T1628;
  wire T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire[7:0] T1634;
  wire[7:0] T1635;
  wire[7:0] T1636;
  reg[7:0] EmitReturnState_3;
  wire T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire T1644;
  wire T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire T1652;
  wire T1653;
  wire[7:0] T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire[7:0] T1663;
  wire[7:0] T1664;
  wire[7:0] T1665;
  reg[7:0] EmitReturnState_2;
  wire T1666;
  wire T1667;
  wire T1668;
  wire T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire T1676;
  wire T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire[7:0] T1683;
  wire T1684;
  wire T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire T1689;
  wire T1690;
  wire T1691;
  wire[7:0] T1692;
  wire[7:0] T1693;
  wire[7:0] T1694;
  reg[7:0] EmitReturnState_1;
  wire T1695;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire T1700;
  wire T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire T1705;
  wire T1706;
  wire T1707;
  wire T1708;
  wire T1709;
  wire T1710;
  wire T1711;
  wire[7:0] T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire T1716;
  wire T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[7:0] T1721;
  wire[7:0] T1722;
  reg[7:0] EmitReturnState_0;
  wire T1723;
  wire T1724;
  wire T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire T1738;
  wire T1739;
  wire[7:0] T1740;
  wire T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire T1745;
  wire T1746;
  wire T1747;
  wire T1748;
  wire[7:0] T1749;
  wire[7:0] T1750;
  wire[7:0] T1751;
  wire[7:0] T1752;
  wire[7:0] T1753;
  wire[7:0] T1754;
  wire[7:0] T1755;
  wire[7:0] T1756;
  wire[7:0] T1757;
  wire[7:0] T1758;
  wire[7:0] T1759;
  wire[7:0] T1760;
  wire[7:0] T1761;
  wire[7:0] T1762;
  wire[7:0] T1763;
  wire[7:0] T1764;
  wire[7:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire T1770;
  wire T1771;
  wire T1772;
  wire T1773;
  wire[7:0] T1774;
  wire[7:0] T1775;
  wire[7:0] T1776;
  reg[7:0] State_4;
  wire T1777;
  wire T1778;
  wire T1779;
  wire T1780;
  wire T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire T1788;
  wire T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire T1796;
  wire T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire T1804;
  wire T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire T1812;
  wire T1813;
  wire[7:0] T1814;
  wire[7:0] T1815;
  wire[7:0] T1816;
  wire[7:0] T1817;
  wire[7:0] T1818;
  wire[7:0] T1819;
  wire[7:0] T1820;
  wire[7:0] T1821;
  wire[7:0] T1822;
  wire[7:0] T1823;
  wire[7:0] T1824;
  wire[7:0] T1825;
  wire[7:0] T1826;
  wire[7:0] T1827;
  wire[7:0] T1828;
  wire[7:0] T1829;
  wire[7:0] T1830;
  wire[7:0] T1831;
  wire[7:0] T1832;
  wire[7:0] T1833;
  wire[7:0] T1834;
  wire[7:0] T1835;
  wire[7:0] T1836;
  wire[7:0] T1837;
  wire[7:0] T1838;
  wire[7:0] T1839;
  wire[7:0] T1840;
  wire[7:0] T1841;
  wire[7:0] T1842;
  wire[7:0] T1843;
  wire[7:0] T1844;
  wire[7:0] T1845;
  wire[7:0] T1846;
  wire[7:0] T1847;
  wire[7:0] T1848;
  wire[7:0] T1849;
  wire[7:0] T1850;
  wire[7:0] T1851;
  wire T1852;
  wire T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire T1859;
  wire[7:0] T1860;
  wire[7:0] T1861;
  wire[7:0] T1862;
  reg[7:0] State_3;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire T1868;
  wire T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire T1884;
  wire T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[7:0] T1900;
  wire[7:0] T1901;
  wire[7:0] T1902;
  wire[7:0] T1903;
  wire[7:0] T1904;
  wire[7:0] T1905;
  wire[7:0] T1906;
  wire[7:0] T1907;
  wire[7:0] T1908;
  wire[7:0] T1909;
  wire[7:0] T1910;
  wire[7:0] T1911;
  wire[7:0] T1912;
  wire[7:0] T1913;
  wire[7:0] T1914;
  wire[7:0] T1915;
  wire[7:0] T1916;
  wire[7:0] T1917;
  wire[7:0] T1918;
  wire[7:0] T1919;
  wire[7:0] T1920;
  wire[7:0] T1921;
  wire[7:0] T1922;
  wire[7:0] T1923;
  wire[7:0] T1924;
  wire[7:0] T1925;
  wire[7:0] T1926;
  wire[7:0] T1927;
  wire[7:0] T1928;
  wire[7:0] T1929;
  wire[7:0] T1930;
  wire[7:0] T1931;
  wire[7:0] T1932;
  wire[7:0] T1933;
  wire[7:0] T1934;
  wire[7:0] T1935;
  wire[7:0] T1936;
  wire[7:0] T1937;
  wire T1938;
  wire T1939;
  wire T1940;
  wire T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire T1945;
  wire[7:0] T1946;
  wire[7:0] T1947;
  wire[7:0] T1948;
  reg[7:0] State_2;
  wire T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire T1955;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire T1972;
  wire T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire T1985;
  wire[7:0] T1986;
  wire[7:0] T1987;
  wire[7:0] T1988;
  wire[7:0] T1989;
  wire[7:0] T1990;
  wire[7:0] T1991;
  wire[7:0] T1992;
  wire[7:0] T1993;
  wire[7:0] T1994;
  wire[7:0] T1995;
  wire[7:0] T1996;
  wire[7:0] T1997;
  wire[7:0] T1998;
  wire[7:0] T1999;
  wire[7:0] T2000;
  wire[7:0] T2001;
  wire[7:0] T2002;
  wire[7:0] T2003;
  wire[7:0] T2004;
  wire[7:0] T2005;
  wire[7:0] T2006;
  wire[7:0] T2007;
  wire[7:0] T2008;
  wire[7:0] T2009;
  wire[7:0] T2010;
  wire[7:0] T2011;
  wire[7:0] T2012;
  wire[7:0] T2013;
  wire[7:0] T2014;
  wire[7:0] T2015;
  wire[7:0] T2016;
  wire[7:0] T2017;
  wire[7:0] T2018;
  wire[7:0] T2019;
  wire[7:0] T2020;
  wire[7:0] T2021;
  wire[7:0] T2022;
  wire[7:0] T2023;
  wire T2024;
  wire T2025;
  wire T2026;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire[7:0] T2032;
  wire[7:0] T2033;
  wire[7:0] T2034;
  reg[7:0] State_1;
  wire T2035;
  wire T2036;
  wire T2037;
  wire T2038;
  wire T2039;
  wire T2040;
  wire T2041;
  wire T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  wire T2051;
  wire T2052;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  wire T2057;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire T2065;
  wire T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire T2070;
  wire T2071;
  wire[7:0] T2072;
  wire[7:0] T2073;
  wire[7:0] T2074;
  wire[7:0] T2075;
  wire[7:0] T2076;
  wire[7:0] T2077;
  wire[7:0] T2078;
  wire[7:0] T2079;
  wire[7:0] T2080;
  wire[7:0] T2081;
  wire[7:0] T2082;
  wire[7:0] T2083;
  wire[7:0] T2084;
  wire[7:0] T2085;
  wire[7:0] T2086;
  wire[7:0] T2087;
  wire[7:0] T2088;
  wire[7:0] T2089;
  wire[7:0] T2090;
  wire[7:0] T2091;
  wire[7:0] T2092;
  wire[7:0] T2093;
  wire[7:0] T2094;
  wire[7:0] T2095;
  wire[7:0] T2096;
  wire[7:0] T2097;
  wire[7:0] T2098;
  wire[7:0] T2099;
  wire[7:0] T2100;
  wire[7:0] T2101;
  wire[7:0] T2102;
  wire[7:0] T2103;
  wire[7:0] T2104;
  wire[7:0] T2105;
  wire[7:0] T2106;
  wire[7:0] T2107;
  wire[7:0] T2108;
  wire[7:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire T2115;
  wire T2116;
  wire T2117;
  wire[7:0] T2118;
  wire[7:0] T2119;
  reg[7:0] State_0;
  wire T2120;
  wire T2121;
  wire T2122;
  wire T2123;
  wire T2124;
  wire T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire T2139;
  wire T2140;
  wire T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire[7:0] T2157;
  wire[7:0] T2158;
  wire[7:0] T2159;
  wire[7:0] T2160;
  wire[7:0] T2161;
  wire[7:0] T2162;
  wire[7:0] T2163;
  wire[7:0] T2164;
  wire[7:0] T2165;
  wire[7:0] T2166;
  wire[7:0] T2167;
  wire[7:0] T2168;
  wire[7:0] T2169;
  wire[7:0] T2170;
  wire[7:0] T2171;
  wire[7:0] T2172;
  wire[7:0] T2173;
  wire[7:0] T2174;
  wire[7:0] T2175;
  wire[7:0] T2176;
  wire[7:0] T2177;
  wire[7:0] T2178;
  wire[7:0] T2179;
  wire[7:0] T2180;
  wire[7:0] T2181;
  wire[7:0] T2182;
  wire[7:0] T2183;
  wire[7:0] T2184;
  wire[7:0] T2185;
  wire[7:0] T2186;
  wire[7:0] T2187;
  wire[7:0] T2188;
  wire[7:0] T2189;
  wire[7:0] T2190;
  wire[7:0] T2191;
  wire[7:0] T2192;
  wire[7:0] T2193;
  wire[7:0] T2194;
  wire T2195;
  wire T2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire T2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  wire T2211;
  wire T2212;
  wire T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  wire T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire T2225;
  wire T2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  wire T2236;
  wire T2237;
  wire T2238;
  wire T2239;
  wire[7:0] T2240;
  wire[7:0] T2241;
  wire[7:0] T2242;
  wire[7:0] T2243;
  wire[7:0] T2244;
  wire[7:0] T2245;
  wire[7:0] T2246;
  wire[7:0] T2247;
  wire[7:0] T2248;
  wire[7:0] T2249;
  wire[7:0] T2250;
  wire[7:0] T2251;
  wire[7:0] T2252;
  wire[7:0] T2253;
  wire[7:0] T2254;
  wire[7:0] T2255;
  wire[7:0] T2256;
  wire[7:0] T2257;
  wire[7:0] T2258;
  wire[7:0] T2259;
  wire[7:0] T2260;
  wire[7:0] T2261;
  wire[7:0] T2262;
  wire[7:0] T2263;
  wire[7:0] T2264;
  wire[7:0] T2265;
  wire[7:0] T2266;
  wire[7:0] T2267;
  wire[7:0] T2268;
  wire[7:0] T2269;
  wire[7:0] T2270;
  wire[7:0] T2271;
  wire[7:0] T2272;
  wire[7:0] T2273;
  wire[7:0] T2274;
  wire[7:0] T2275;
  wire[7:0] T2276;
  wire[7:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire T2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire T2289;
  wire[3:0] T2290;
  wire T2291;
  reg[0:0] subStateTh_5;
  wire T2292;
  wire T2293;
  wire T2294;
  wire[3:0] T2295;
  wire T2296;
  wire T2297;
  wire T2298;
  wire T2299;
  wire T2300;
  wire T2301;
  wire[3:0] T2302;
  wire T2303;
  reg[0:0] subStateTh_4;
  wire T2304;
  wire T2305;
  wire T2306;
  wire[3:0] T2307;
  wire T2308;
  wire T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire T2313;
  wire[3:0] T2314;
  wire T2315;
  reg[0:0] subStateTh_3;
  wire T2316;
  wire T2317;
  wire T2318;
  wire[3:0] T2319;
  wire T2320;
  wire T2321;
  wire T2322;
  wire T2323;
  wire T2324;
  wire T2325;
  wire[3:0] T2326;
  wire T2327;
  reg[0:0] subStateTh_2;
  wire T2328;
  wire T2329;
  wire T2330;
  wire[3:0] T2331;
  wire T2332;
  wire T2333;
  wire T2334;
  wire T2335;
  wire T2336;
  wire T2337;
  wire[3:0] T2338;
  wire T2339;
  reg[0:0] subStateTh_1;
  wire T2340;
  wire T2341;
  wire T2342;
  wire[3:0] T2343;
  wire T2344;
  wire T2345;
  wire T2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire[3:0] T2350;
  wire T2351;
  reg[0:0] subStateTh_0;
  wire T2352;
  wire T2353;
  wire T2354;
  wire[3:0] T2355;
  wire T2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  wire T2361;
  wire[3:0] T2362;
  wire T2363;
  wire[7:0] T2364;
  wire[7:0] T2365;
  wire[7:0] T2366;
  wire[7:0] T2367;
  wire[7:0] T2368;
  wire[7:0] T2369;
  wire[7:0] T2370;
  wire[7:0] T2371;
  wire[7:0] T2372;
  wire[7:0] T2373;
  wire[7:0] T2374;
  wire[7:0] T2375;
  wire[7:0] T2376;
  wire[7:0] T2377;
  wire[7:0] T2378;
  wire[7:0] T2379;
  wire[7:0] T2380;
  wire[7:0] T2381;
  wire[7:0] T2382;
  wire[7:0] T2383;
  wire T2384;
  wire T2385;
  wire T2386;
  wire T2387;
  wire T2388;
  reg[0:0] dramBank7_valid_received_7;
  wire T2389;
  wire T2390;
  wire T2391;
  wire T2392;
  wire[9:0] T2393;
  wire[9:0] dramBank7Port_rep_tag;
  wire[9:0] dramBank7Port_req_tag;
  wire[9:0] T2394;
  wire dramBank7Port_rep_valid;
  wire T2395;
  wire T2396;
  wire[4:0] T2397;
  wire T2398;
  wire T2399;
  reg[0:0] dramBank7_valid_received_6;
  wire T2400;
  wire T2401;
  wire T2402;
  wire T2403;
  wire[9:0] T2404;
  wire T2405;
  wire T2406;
  wire[4:0] T2407;
  wire T2408;
  wire T2409;
  reg[0:0] dramBank7_valid_received_5;
  wire T2410;
  wire T2411;
  wire T2412;
  wire T2413;
  wire[9:0] T2414;
  wire T2415;
  wire T2416;
  wire[4:0] T2417;
  wire T2418;
  wire T2419;
  reg[0:0] dramBank7_valid_received_4;
  wire T2420;
  wire T2421;
  wire T2422;
  wire T2423;
  wire[9:0] T2424;
  wire T2425;
  wire T2426;
  wire[4:0] T2427;
  wire T2428;
  wire T2429;
  reg[0:0] dramBank7_valid_received_3;
  wire T2430;
  wire T2431;
  wire T2432;
  wire T2433;
  wire[9:0] T2434;
  wire T2435;
  wire T2436;
  wire[4:0] T2437;
  wire T2438;
  wire T2439;
  reg[0:0] dramBank7_valid_received_2;
  wire T2440;
  wire T2441;
  wire T2442;
  wire T2443;
  wire[9:0] T2444;
  wire T2445;
  wire T2446;
  wire[4:0] T2447;
  wire T2448;
  wire T2449;
  reg[0:0] dramBank7_valid_received_1;
  wire T2450;
  wire T2451;
  wire T2452;
  wire T2453;
  wire[9:0] T2454;
  wire T2455;
  wire T2456;
  wire[4:0] T2457;
  wire T2458;
  reg[0:0] dramBank7_valid_received_0;
  wire T2459;
  wire T2460;
  wire T2461;
  wire T2462;
  wire[9:0] T2463;
  wire T2464;
  wire T2465;
  wire[4:0] T2466;
  wire T2467;
  wire T2468;
  wire[4:0] T2469;
  wire T2470;
  wire T2471;
  wire[4:0] T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  wire[9:0] T2476;
  wire T2477;
  wire T2478;
  wire T2479;
  reg[0:0] dramBank6PortHadValidRequest_7;
  wire T2480;
  wire T2481;
  wire T2482;
  wire T2483;
  wire[4:0] T2484;
  wire T2485;
  wire T2486;
  wire[4:0] T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  wire[9:0] T2491;
  wire T2492;
  wire T2493;
  wire T2494;
  reg[0:0] dramBank5PortHadValidRequest_7;
  wire T2495;
  wire T2496;
  wire T2497;
  wire T2498;
  wire[4:0] T2499;
  wire T2500;
  wire T2501;
  wire[4:0] T2502;
  wire T2503;
  wire T2504;
  wire T2505;
  wire[9:0] T2506;
  wire T2507;
  wire T2508;
  wire T2509;
  reg[0:0] dramBank4PortHadValidRequest_7;
  wire T2510;
  wire T2511;
  wire T2512;
  wire T2513;
  wire[4:0] T2514;
  wire T2515;
  wire T2516;
  wire[4:0] T2517;
  wire T2518;
  wire T2519;
  wire T2520;
  wire[9:0] T2521;
  wire T2522;
  wire T2523;
  wire T2524;
  reg[0:0] dramBank3PortHadValidRequest_7;
  wire T2525;
  wire T2526;
  wire T2527;
  wire T2528;
  wire[4:0] T2529;
  wire T2530;
  wire T2531;
  wire[4:0] T2532;
  wire T2533;
  wire T2534;
  wire T2535;
  wire[9:0] T2536;
  wire T2537;
  wire T2538;
  wire T2539;
  reg[0:0] dramBank2PortHadValidRequest_7;
  wire T2540;
  wire T2541;
  wire T2542;
  wire T2543;
  wire[4:0] T2544;
  wire T2545;
  wire T2546;
  wire[4:0] T2547;
  wire T2548;
  wire T2549;
  wire T2550;
  wire[9:0] T2551;
  wire T2552;
  wire T2553;
  wire T2554;
  reg[0:0] dramBank1PortHadValidRequest_7;
  wire T2555;
  wire T2556;
  wire T2557;
  wire T2558;
  wire[4:0] T2559;
  wire T2560;
  wire T2561;
  wire[4:0] T2562;
  wire T2563;
  wire T2564;
  wire T2565;
  wire[9:0] T2566;
  wire T2567;
  wire T2568;
  reg[0:0] dramBank0PortHadValidRequest_7;
  wire T2569;
  wire T2570;
  wire T2571;
  wire T2572;
  wire[4:0] T2573;
  wire T2574;
  wire T2575;
  wire[4:0] T2576;
  wire T2577;
  wire T2578;
  wire T2579;
  wire[9:0] T2580;
  wire T2581;
  wire T2582;
  wire AllOffloadsValid_6;
  wire T2583;
  wire T2584;
  wire T2585;
  reg[0:0] dramBank7PortHadValidRequest_6;
  wire T2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire[4:0] T2590;
  wire T2591;
  wire T2592;
  wire[4:0] T2593;
  wire T2594;
  wire T2595;
  wire T2596;
  wire[9:0] T2597;
  wire T2598;
  wire T2599;
  wire T2600;
  reg[0:0] dramBank6PortHadValidRequest_6;
  wire T2601;
  wire T2602;
  wire T2603;
  wire T2604;
  wire[4:0] T2605;
  wire T2606;
  wire T2607;
  wire[4:0] T2608;
  wire T2609;
  wire T2610;
  wire T2611;
  wire[9:0] T2612;
  wire T2613;
  wire T2614;
  wire T2615;
  reg[0:0] dramBank5PortHadValidRequest_6;
  wire T2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire[4:0] T2620;
  wire T2621;
  wire T2622;
  wire[4:0] T2623;
  wire T2624;
  wire T2625;
  wire T2626;
  wire[9:0] T2627;
  wire T2628;
  wire T2629;
  wire T2630;
  reg[0:0] dramBank4PortHadValidRequest_6;
  wire T2631;
  wire T2632;
  wire T2633;
  wire T2634;
  wire[4:0] T2635;
  wire T2636;
  wire T2637;
  wire[4:0] T2638;
  wire T2639;
  wire T2640;
  wire T2641;
  wire[9:0] T2642;
  wire T2643;
  wire T2644;
  wire T2645;
  reg[0:0] dramBank3PortHadValidRequest_6;
  wire T2646;
  wire T2647;
  wire T2648;
  wire T2649;
  wire[4:0] T2650;
  wire T2651;
  wire T2652;
  wire[4:0] T2653;
  wire T2654;
  wire T2655;
  wire T2656;
  wire[9:0] T2657;
  wire T2658;
  wire T2659;
  wire T2660;
  reg[0:0] dramBank2PortHadValidRequest_6;
  wire T2661;
  wire T2662;
  wire T2663;
  wire T2664;
  wire[4:0] T2665;
  wire T2666;
  wire T2667;
  wire[4:0] T2668;
  wire T2669;
  wire T2670;
  wire T2671;
  wire[9:0] T2672;
  wire T2673;
  wire T2674;
  wire T2675;
  reg[0:0] dramBank1PortHadValidRequest_6;
  wire T2676;
  wire T2677;
  wire T2678;
  wire T2679;
  wire[4:0] T2680;
  wire T2681;
  wire T2682;
  wire[4:0] T2683;
  wire T2684;
  wire T2685;
  wire T2686;
  wire[9:0] T2687;
  wire T2688;
  wire T2689;
  reg[0:0] dramBank0PortHadValidRequest_6;
  wire T2690;
  wire T2691;
  wire T2692;
  wire T2693;
  wire[4:0] T2694;
  wire T2695;
  wire T2696;
  wire[4:0] T2697;
  wire T2698;
  wire T2699;
  wire T2700;
  wire[9:0] T2701;
  wire T2702;
  wire T2703;
  wire AllOffloadsValid_5;
  wire T2704;
  wire T2705;
  wire T2706;
  reg[0:0] dramBank7PortHadValidRequest_5;
  wire T2707;
  wire T2708;
  wire T2709;
  wire T2710;
  wire[4:0] T2711;
  wire T2712;
  wire T2713;
  wire[4:0] T2714;
  wire T2715;
  wire T2716;
  wire T2717;
  wire[9:0] T2718;
  wire T2719;
  wire T2720;
  wire T2721;
  reg[0:0] dramBank6PortHadValidRequest_5;
  wire T2722;
  wire T2723;
  wire T2724;
  wire T2725;
  wire[4:0] T2726;
  wire T2727;
  wire T2728;
  wire[4:0] T2729;
  wire T2730;
  wire T2731;
  wire T2732;
  wire[9:0] T2733;
  wire T2734;
  wire T2735;
  wire T2736;
  reg[0:0] dramBank5PortHadValidRequest_5;
  wire T2737;
  wire T2738;
  wire T2739;
  wire T2740;
  wire[4:0] T2741;
  wire T2742;
  wire T2743;
  wire[4:0] T2744;
  wire T2745;
  wire T2746;
  wire T2747;
  wire[9:0] T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  reg[0:0] dramBank4PortHadValidRequest_5;
  wire T2752;
  wire T2753;
  wire T2754;
  wire T2755;
  wire[4:0] T2756;
  wire T2757;
  wire T2758;
  wire[4:0] T2759;
  wire T2760;
  wire T2761;
  wire T2762;
  wire[9:0] T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  reg[0:0] dramBank3PortHadValidRequest_5;
  wire T2767;
  wire T2768;
  wire T2769;
  wire T2770;
  wire[4:0] T2771;
  wire T2772;
  wire T2773;
  wire[4:0] T2774;
  wire T2775;
  wire T2776;
  wire T2777;
  wire[9:0] T2778;
  wire T2779;
  wire T2780;
  wire T2781;
  reg[0:0] dramBank2PortHadValidRequest_5;
  wire T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  wire[4:0] T2786;
  wire T2787;
  wire T2788;
  wire[4:0] T2789;
  wire T2790;
  wire T2791;
  wire T2792;
  wire[9:0] T2793;
  wire T2794;
  wire T2795;
  wire T2796;
  reg[0:0] dramBank1PortHadValidRequest_5;
  wire T2797;
  wire T2798;
  wire T2799;
  wire T2800;
  wire[4:0] T2801;
  wire T2802;
  wire T2803;
  wire[4:0] T2804;
  wire T2805;
  wire T2806;
  wire T2807;
  wire[9:0] T2808;
  wire T2809;
  wire T2810;
  reg[0:0] dramBank0PortHadValidRequest_5;
  wire T2811;
  wire T2812;
  wire T2813;
  wire T2814;
  wire[4:0] T2815;
  wire T2816;
  wire T2817;
  wire[4:0] T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire[9:0] T2822;
  wire T2823;
  wire T2824;
  wire AllOffloadsValid_4;
  wire T2825;
  wire T2826;
  wire T2827;
  reg[0:0] dramBank7PortHadValidRequest_4;
  wire T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire[4:0] T2832;
  wire T2833;
  wire T2834;
  wire[4:0] T2835;
  wire T2836;
  wire T2837;
  wire T2838;
  wire[9:0] T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  reg[0:0] dramBank6PortHadValidRequest_4;
  wire T2843;
  wire T2844;
  wire T2845;
  wire T2846;
  wire[4:0] T2847;
  wire T2848;
  wire T2849;
  wire[4:0] T2850;
  wire T2851;
  wire T2852;
  wire T2853;
  wire[9:0] T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  reg[0:0] dramBank5PortHadValidRequest_4;
  wire T2858;
  wire T2859;
  wire T2860;
  wire T2861;
  wire[4:0] T2862;
  wire T2863;
  wire T2864;
  wire[4:0] T2865;
  wire T2866;
  wire T2867;
  wire T2868;
  wire[9:0] T2869;
  wire T2870;
  wire T2871;
  wire T2872;
  reg[0:0] dramBank4PortHadValidRequest_4;
  wire T2873;
  wire T2874;
  wire T2875;
  wire T2876;
  wire[4:0] T2877;
  wire T2878;
  wire T2879;
  wire[4:0] T2880;
  wire T2881;
  wire T2882;
  wire T2883;
  wire[9:0] T2884;
  wire T2885;
  wire T2886;
  wire T2887;
  reg[0:0] dramBank3PortHadValidRequest_4;
  wire T2888;
  wire T2889;
  wire T2890;
  wire T2891;
  wire[4:0] T2892;
  wire T2893;
  wire T2894;
  wire[4:0] T2895;
  wire T2896;
  wire T2897;
  wire T2898;
  wire[9:0] T2899;
  wire T2900;
  wire T2901;
  wire T2902;
  reg[0:0] dramBank2PortHadValidRequest_4;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire[4:0] T2907;
  wire T2908;
  wire T2909;
  wire[4:0] T2910;
  wire T2911;
  wire T2912;
  wire T2913;
  wire[9:0] T2914;
  wire T2915;
  wire T2916;
  wire T2917;
  reg[0:0] dramBank1PortHadValidRequest_4;
  wire T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire[4:0] T2922;
  wire T2923;
  wire T2924;
  wire[4:0] T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire[9:0] T2929;
  wire T2930;
  wire T2931;
  reg[0:0] dramBank0PortHadValidRequest_4;
  wire T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire[4:0] T2936;
  wire T2937;
  wire T2938;
  wire[4:0] T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire[9:0] T2943;
  wire T2944;
  wire T2945;
  wire AllOffloadsValid_3;
  wire T2946;
  wire T2947;
  wire T2948;
  reg[0:0] dramBank7PortHadValidRequest_3;
  wire T2949;
  wire T2950;
  wire T2951;
  wire T2952;
  wire[4:0] T2953;
  wire T2954;
  wire T2955;
  wire[4:0] T2956;
  wire T2957;
  wire T2958;
  wire T2959;
  wire[9:0] T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  reg[0:0] dramBank6PortHadValidRequest_3;
  wire T2964;
  wire T2965;
  wire T2966;
  wire T2967;
  wire[4:0] T2968;
  wire T2969;
  wire T2970;
  wire[4:0] T2971;
  wire T2972;
  wire T2973;
  wire T2974;
  wire[9:0] T2975;
  wire T2976;
  wire T2977;
  wire T2978;
  reg[0:0] dramBank5PortHadValidRequest_3;
  wire T2979;
  wire T2980;
  wire T2981;
  wire T2982;
  wire[4:0] T2983;
  wire T2984;
  wire T2985;
  wire[4:0] T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire[9:0] T2990;
  wire T2991;
  wire T2992;
  wire T2993;
  reg[0:0] dramBank4PortHadValidRequest_3;
  wire T2994;
  wire T2995;
  wire T2996;
  wire T2997;
  wire[4:0] T2998;
  wire T2999;
  wire T3000;
  wire[4:0] T3001;
  wire T3002;
  wire T3003;
  wire T3004;
  wire[9:0] T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  reg[0:0] dramBank3PortHadValidRequest_3;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire[4:0] T3013;
  wire T3014;
  wire T3015;
  wire[4:0] T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire[9:0] T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  reg[0:0] dramBank2PortHadValidRequest_3;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire[4:0] T3028;
  wire T3029;
  wire T3030;
  wire[4:0] T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire[9:0] T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  reg[0:0] dramBank1PortHadValidRequest_3;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire[4:0] T3043;
  wire T3044;
  wire T3045;
  wire[4:0] T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire[9:0] T3050;
  wire T3051;
  wire T3052;
  reg[0:0] dramBank0PortHadValidRequest_3;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire[4:0] T3057;
  wire T3058;
  wire T3059;
  wire[4:0] T3060;
  wire T3061;
  wire T3062;
  wire T3063;
  wire[9:0] T3064;
  wire T3065;
  wire T3066;
  wire AllOffloadsValid_2;
  wire T3067;
  wire T3068;
  wire T3069;
  reg[0:0] dramBank7PortHadValidRequest_2;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire[4:0] T3074;
  wire T3075;
  wire T3076;
  wire[4:0] T3077;
  wire T3078;
  wire T3079;
  wire T3080;
  wire[9:0] T3081;
  wire T3082;
  wire T3083;
  wire T3084;
  reg[0:0] dramBank6PortHadValidRequest_2;
  wire T3085;
  wire T3086;
  wire T3087;
  wire T3088;
  wire[4:0] T3089;
  wire T3090;
  wire T3091;
  wire[4:0] T3092;
  wire T3093;
  wire T3094;
  wire T3095;
  wire[9:0] T3096;
  wire T3097;
  wire T3098;
  wire T3099;
  reg[0:0] dramBank5PortHadValidRequest_2;
  wire T3100;
  wire T3101;
  wire T3102;
  wire T3103;
  wire[4:0] T3104;
  wire T3105;
  wire T3106;
  wire[4:0] T3107;
  wire T3108;
  wire T3109;
  wire T3110;
  wire[9:0] T3111;
  wire T3112;
  wire T3113;
  wire T3114;
  reg[0:0] dramBank4PortHadValidRequest_2;
  wire T3115;
  wire T3116;
  wire T3117;
  wire T3118;
  wire[4:0] T3119;
  wire T3120;
  wire T3121;
  wire[4:0] T3122;
  wire T3123;
  wire T3124;
  wire T3125;
  wire[9:0] T3126;
  wire T3127;
  wire T3128;
  wire T3129;
  reg[0:0] dramBank3PortHadValidRequest_2;
  wire T3130;
  wire T3131;
  wire T3132;
  wire T3133;
  wire[4:0] T3134;
  wire T3135;
  wire T3136;
  wire[4:0] T3137;
  wire T3138;
  wire T3139;
  wire T3140;
  wire[9:0] T3141;
  wire T3142;
  wire T3143;
  wire T3144;
  reg[0:0] dramBank2PortHadValidRequest_2;
  wire T3145;
  wire T3146;
  wire T3147;
  wire T3148;
  wire[4:0] T3149;
  wire T3150;
  wire T3151;
  wire[4:0] T3152;
  wire T3153;
  wire T3154;
  wire T3155;
  wire[9:0] T3156;
  wire T3157;
  wire T3158;
  wire T3159;
  reg[0:0] dramBank1PortHadValidRequest_2;
  wire T3160;
  wire T3161;
  wire T3162;
  wire T3163;
  wire[4:0] T3164;
  wire T3165;
  wire T3166;
  wire[4:0] T3167;
  wire T3168;
  wire T3169;
  wire T3170;
  wire[9:0] T3171;
  wire T3172;
  wire T3173;
  reg[0:0] dramBank0PortHadValidRequest_2;
  wire T3174;
  wire T3175;
  wire T3176;
  wire T3177;
  wire[4:0] T3178;
  wire T3179;
  wire T3180;
  wire[4:0] T3181;
  wire T3182;
  wire T3183;
  wire T3184;
  wire[9:0] T3185;
  wire T3186;
  wire T3187;
  wire AllOffloadsValid_1;
  wire T3188;
  wire T3189;
  wire T3190;
  reg[0:0] dramBank7PortHadValidRequest_1;
  wire T3191;
  wire T3192;
  wire T3193;
  wire T3194;
  wire[4:0] T3195;
  wire T3196;
  wire T3197;
  wire[4:0] T3198;
  wire T3199;
  wire T3200;
  wire T3201;
  wire[9:0] T3202;
  wire T3203;
  wire T3204;
  wire T3205;
  reg[0:0] dramBank6PortHadValidRequest_1;
  wire T3206;
  wire T3207;
  wire T3208;
  wire T3209;
  wire[4:0] T3210;
  wire T3211;
  wire T3212;
  wire[4:0] T3213;
  wire T3214;
  wire T3215;
  wire T3216;
  wire[9:0] T3217;
  wire T3218;
  wire T3219;
  wire T3220;
  reg[0:0] dramBank5PortHadValidRequest_1;
  wire T3221;
  wire T3222;
  wire T3223;
  wire T3224;
  wire[4:0] T3225;
  wire T3226;
  wire T3227;
  wire[4:0] T3228;
  wire T3229;
  wire T3230;
  wire T3231;
  wire[9:0] T3232;
  wire T3233;
  wire T3234;
  wire T3235;
  reg[0:0] dramBank4PortHadValidRequest_1;
  wire T3236;
  wire T3237;
  wire T3238;
  wire T3239;
  wire[4:0] T3240;
  wire T3241;
  wire T3242;
  wire[4:0] T3243;
  wire T3244;
  wire T3245;
  wire T3246;
  wire[9:0] T3247;
  wire T3248;
  wire T3249;
  wire T3250;
  reg[0:0] dramBank3PortHadValidRequest_1;
  wire T3251;
  wire T3252;
  wire T3253;
  wire T3254;
  wire[4:0] T3255;
  wire T3256;
  wire T3257;
  wire[4:0] T3258;
  wire T3259;
  wire T3260;
  wire T3261;
  wire[9:0] T3262;
  wire T3263;
  wire T3264;
  wire T3265;
  reg[0:0] dramBank2PortHadValidRequest_1;
  wire T3266;
  wire T3267;
  wire T3268;
  wire T3269;
  wire[4:0] T3270;
  wire T3271;
  wire T3272;
  wire[4:0] T3273;
  wire T3274;
  wire T3275;
  wire T3276;
  wire[9:0] T3277;
  wire T3278;
  wire T3279;
  wire T3280;
  reg[0:0] dramBank1PortHadValidRequest_1;
  wire T3281;
  wire T3282;
  wire T3283;
  wire T3284;
  wire[4:0] T3285;
  wire T3286;
  wire T3287;
  wire[4:0] T3288;
  wire T3289;
  wire T3290;
  wire T3291;
  wire[9:0] T3292;
  wire T3293;
  wire T3294;
  reg[0:0] dramBank0PortHadValidRequest_1;
  wire T3295;
  wire T3296;
  wire T3297;
  wire T3298;
  wire[4:0] T3299;
  wire T3300;
  wire T3301;
  wire[4:0] T3302;
  wire T3303;
  wire T3304;
  wire T3305;
  wire[9:0] T3306;
  wire T3307;
  wire T3308;
  wire AllOffloadsValid_0;
  wire T3309;
  wire T3310;
  wire T3311;
  reg[0:0] dramBank7PortHadValidRequest_0;
  wire T3312;
  wire T3313;
  wire T3314;
  wire T3315;
  wire[4:0] T3316;
  wire T3317;
  wire T3318;
  wire[4:0] T3319;
  wire T3320;
  wire T3321;
  wire T3322;
  wire[9:0] T3323;
  wire T3324;
  wire T3325;
  wire T3326;
  reg[0:0] dramBank6PortHadValidRequest_0;
  wire T3327;
  wire T3328;
  wire T3329;
  wire T3330;
  wire[4:0] T3331;
  wire T3332;
  wire T3333;
  wire[4:0] T3334;
  wire T3335;
  wire T3336;
  wire T3337;
  wire[9:0] T3338;
  wire T3339;
  wire T3340;
  wire T3341;
  reg[0:0] dramBank5PortHadValidRequest_0;
  wire T3342;
  wire T3343;
  wire T3344;
  wire T3345;
  wire[4:0] T3346;
  wire T3347;
  wire T3348;
  wire[4:0] T3349;
  wire T3350;
  wire T3351;
  wire T3352;
  wire[9:0] T3353;
  wire T3354;
  wire T3355;
  wire T3356;
  reg[0:0] dramBank4PortHadValidRequest_0;
  wire T3357;
  wire T3358;
  wire T3359;
  wire T3360;
  wire[4:0] T3361;
  wire T3362;
  wire T3363;
  wire[4:0] T3364;
  wire T3365;
  wire T3366;
  wire T3367;
  wire[9:0] T3368;
  wire T3369;
  wire T3370;
  wire T3371;
  reg[0:0] dramBank3PortHadValidRequest_0;
  wire T3372;
  wire T3373;
  wire T3374;
  wire T3375;
  wire[4:0] T3376;
  wire T3377;
  wire T3378;
  wire[4:0] T3379;
  wire T3380;
  wire T3381;
  wire T3382;
  wire[9:0] T3383;
  wire T3384;
  wire T3385;
  wire T3386;
  reg[0:0] dramBank2PortHadValidRequest_0;
  wire T3387;
  wire T3388;
  wire T3389;
  wire T3390;
  wire[4:0] T3391;
  wire T3392;
  wire T3393;
  wire[4:0] T3394;
  wire T3395;
  wire T3396;
  wire T3397;
  wire[9:0] T3398;
  wire T3399;
  wire T3400;
  wire T3401;
  reg[0:0] dramBank1PortHadValidRequest_0;
  wire T3402;
  wire T3403;
  wire T3404;
  wire T3405;
  wire[4:0] T3406;
  wire T3407;
  wire T3408;
  wire[4:0] T3409;
  wire T3410;
  wire T3411;
  wire T3412;
  wire[9:0] T3413;
  wire T3414;
  wire T3415;
  reg[0:0] dramBank0PortHadValidRequest_0;
  wire T3416;
  wire T3417;
  wire T3418;
  wire T3419;
  wire[4:0] T3420;
  wire T3421;
  wire T3422;
  wire[4:0] T3423;
  wire T3424;
  wire T3425;
  wire T3426;
  wire[9:0] T3427;
  wire T3428;
  wire T3429;
  wire T3430;
  wire T3431;
  wire T3432;
  wire T3433;
  wire T3434;
  wire T3435;
  wire T3436;
  wire T3437;
  wire T3438;
  wire T3439;
  wire T3440;
  wire T3441;
  wire T3442;
  wire T3443;
  wire T3444;
  wire T3445;
  wire T3446;
  wire T3447;
  wire T3448;
  wire T3449;
  wire T3450;
  wire T3451;
  wire T3452;
  wire T3453;
  wire T3454;
  wire T3455;
  wire T3456;
  wire T3457;
  wire T3458;
  wire T3459;
  wire T3460;
  wire T3461;
  wire T3462;
  wire T3463;
  wire T3464;
  wire T3465;
  wire[7:0] T3466;
  wire[7:0] T3467;
  wire[7:0] T3468;
  wire[7:0] T3469;
  wire[7:0] T3470;
  wire[7:0] T3471;
  wire[7:0] T3472;
  wire[7:0] T3473;
  wire[7:0] T3474;
  wire[7:0] T3475;
  wire[7:0] T3476;
  wire[7:0] T3477;
  wire[7:0] T3478;
  wire[7:0] T3479;
  wire[7:0] T3480;
  wire[7:0] T3481;
  wire[7:0] T3482;
  wire[7:0] T3483;
  wire[7:0] T3484;
  wire[7:0] T3485;
  wire[7:0] T3486;
  wire[7:0] T3487;
  wire[7:0] T3488;
  wire[7:0] T3489;
  wire[7:0] T3490;
  wire[7:0] T3491;
  wire[7:0] T3492;
  wire[7:0] T3493;
  wire[7:0] T3494;
  wire[7:0] T3495;
  wire[7:0] T3496;
  wire[7:0] T3497;
  wire[7:0] T3498;
  wire[7:0] T3499;
  wire[7:0] T3500;
  wire[7:0] T3501;
  wire[7:0] T3502;
  wire[7:0] T3503;
  wire T3504;
  wire T3505;
  wire T3506;
  wire T3507;
  wire T3508;
  wire T3509;
  wire T3510;
  wire T3511;
  wire T3512;
  wire T3513;
  wire T3514;
  wire T3515;
  wire T3516;
  wire T3517;
  wire T3518;
  wire T3519;
  wire T3520;
  wire T3521;
  wire T3522;
  wire T3523;
  wire T3524;
  wire T3525;
  wire T3526;
  wire T3527;
  wire T3528;
  wire T3529;
  wire T3530;
  wire T3531;
  wire T3532;
  wire T3533;
  wire T3534;
  wire[9:0] T3535;
  wire[9:0] T3536;
  wire[9:0] T3537;
  reg[9:0] inputTag_7;
  wire[9:0] T3538;
  wire[9:0] T3539;
  wire[9:0] T3540;
  wire[9:0] T3541;
  reg[9:0] inputTag_6;
  wire[9:0] T3542;
  wire[9:0] T3543;
  wire[9:0] T3544;
  wire[9:0] T3545;
  reg[9:0] inputTag_5;
  wire[9:0] T3546;
  wire[9:0] T3547;
  wire[9:0] T3548;
  wire[9:0] T3549;
  reg[9:0] inputTag_4;
  wire[9:0] T3550;
  wire[9:0] T3551;
  wire[9:0] T3552;
  wire[9:0] T3553;
  reg[9:0] inputTag_3;
  wire[9:0] T3554;
  wire[9:0] T3555;
  wire[9:0] T3556;
  wire[9:0] T3557;
  reg[9:0] inputTag_2;
  wire[9:0] T3558;
  wire[9:0] T3559;
  wire[9:0] T3560;
  wire[9:0] T3561;
  reg[9:0] inputTag_1;
  wire[9:0] T3562;
  wire[9:0] T3563;
  wire[9:0] T3564;
  reg[9:0] inputTag_0;
  wire[9:0] T3565;
  wire T3566;
  wire T3567;
  wire T3568;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T1 = T3512 && T2;
  assign T2 = State_7 == 8'h0/* 0*/;
  assign T3 = T3430 || T4;
  assign T4 = T765 && T5;
  assign T5 = T6[3'h7/* 7*/];
  assign T6 = T7[3'h7/* 7*/:1'h0/* 0*/];
  assign T7 = 8'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T2581 && AllOffloadsValid_7;
  assign AllOffloadsValid_7 = T9;
  assign T9 = T2477 && T10;
  assign T10 = T2473 || T11;
  assign T11 = ! dramBank7PortHadValidRequest_7;
  assign T12 = T2470 && T13;
  assign T13 = dramBank7PortHadValidRequest_7 || T14;
  assign T14 = T2468 && dramBank7Port_req_valid;
  assign dramBank7Port_req_valid = T15;
  assign T15 = T2385 && T16;
  assign T16 = T2384 && T17;
  assign T17 = T19 == T18;
  assign T18 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T19 = T2364 | T20;
  assign T20 = State_7 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23[3'h7/* 7*/];
  assign T23 = T24[3'h7/* 7*/:1'h0/* 0*/];
  assign T24 = 8'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_7 == 1'h0/* 0*/;
  assign T26 = T30 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_7;
  assign T28 = T29 == vThreadEncoder_io_chosen;
  assign T29 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T30 = T32 && T31;
  assign T31 = State_7 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_7 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = T36 == rThreadEncoder_io_chosen;
  assign T36 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign AllOffloadsReady = T37;
  assign T37 = T49 && T38;
  assign T38 = T45 || T39;
  assign T39 = T41 && T40;
  assign T40 = ! dramBank7Port_req_valid;
  assign T41 = ! dramBank7PortHadReadyRequest;
  assign T42 = T44 && T43;
  assign T43 = dramBank7PortHadReadyRequest || dramBank7Port_req_valid;
  assign T44 = ! AllOffloadsReady;
  assign T45 = dramBank7Port_req_ready || dramBank7_ready_received;
  assign T46 = T48 && T47;
  assign T47 = dramBank7_ready_received || dramBank7Port_req_ready;
  assign dramBank7Port_req_ready = mainOff_dramBank7_req_ready;
  assign mainOff_dramBank7_rep_ready = dramBank7Port_rep_ready;
  assign dramBank7Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank7_req_valid = dramBank7Port_req_valid;
  assign T48 = ! AllOffloadsReady;
  assign T49 = T156 && T50;
  assign T50 = T152 || T51;
  assign T51 = T148 && T52;
  assign T52 = ! dramBank6Port_req_valid;
  assign dramBank6Port_req_valid = T53;
  assign T53 = T58 && T54;
  assign T54 = T57 && T55;
  assign T55 = T19 == T56;
  assign T56 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T57 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T58 = T147 && T59;
  assign T59 = ! T60;
  assign T60 = T71 | T61;
  assign T61 = dramBank6_valid_received_7 & T22;
  assign T62 = T68 && T63;
  assign T63 = dramBank6_valid_received_7 || T64;
  assign T64 = dramBank6Port_rep_valid && T65;
  assign T65 = dramBank6Port_rep_tag == T66;
  assign T66 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank6Port_rep_tag = mainOff_dramBank6_rep_tag;
  assign mainOff_dramBank6_rep_ready = dramBank6Port_rep_ready;
  assign dramBank6Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank6_req_valid = dramBank6Port_req_valid;
  assign mainOff_dramBank6_req_tag = dramBank6Port_req_tag;
  assign dramBank6Port_req_tag = T67;
  assign T67 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank6Port_rep_valid = mainOff_dramBank6_rep_valid;
  assign T68 = ! T69;
  assign T69 = T70 == 5'h7/* 7*/;
  assign T70 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T71 = T82 | T72;
  assign T72 = dramBank6_valid_received_6 & T73;
  assign T73 = T23[3'h6/* 6*/];
  assign T74 = T79 && T75;
  assign T75 = dramBank6_valid_received_6 || T76;
  assign T76 = dramBank6Port_rep_valid && T77;
  assign T77 = dramBank6Port_rep_tag == T78;
  assign T78 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T79 = ! T80;
  assign T80 = T81 == 5'h6/* 6*/;
  assign T81 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T82 = T93 | T83;
  assign T83 = dramBank6_valid_received_5 & T84;
  assign T84 = T23[3'h5/* 5*/];
  assign T85 = T90 && T86;
  assign T86 = dramBank6_valid_received_5 || T87;
  assign T87 = dramBank6Port_rep_valid && T88;
  assign T88 = dramBank6Port_rep_tag == T89;
  assign T89 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T90 = ! T91;
  assign T91 = T92 == 5'h5/* 5*/;
  assign T92 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T93 = T104 | T94;
  assign T94 = dramBank6_valid_received_4 & T95;
  assign T95 = T23[3'h4/* 4*/];
  assign T96 = T101 && T97;
  assign T97 = dramBank6_valid_received_4 || T98;
  assign T98 = dramBank6Port_rep_valid && T99;
  assign T99 = dramBank6Port_rep_tag == T100;
  assign T100 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T101 = ! T102;
  assign T102 = T103 == 5'h4/* 4*/;
  assign T103 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T104 = T115 | T105;
  assign T105 = dramBank6_valid_received_3 & T106;
  assign T106 = T23[2'h3/* 3*/];
  assign T107 = T112 && T108;
  assign T108 = dramBank6_valid_received_3 || T109;
  assign T109 = dramBank6Port_rep_valid && T110;
  assign T110 = dramBank6Port_rep_tag == T111;
  assign T111 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T112 = ! T113;
  assign T113 = T114 == 5'h3/* 3*/;
  assign T114 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T115 = T126 | T116;
  assign T116 = dramBank6_valid_received_2 & T117;
  assign T117 = T23[2'h2/* 2*/];
  assign T118 = T123 && T119;
  assign T119 = dramBank6_valid_received_2 || T120;
  assign T120 = dramBank6Port_rep_valid && T121;
  assign T121 = dramBank6Port_rep_tag == T122;
  assign T122 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T123 = ! T124;
  assign T124 = T125 == 5'h2/* 2*/;
  assign T125 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T126 = T137 | T127;
  assign T127 = dramBank6_valid_received_1 & T128;
  assign T128 = T23[1'h1/* 1*/];
  assign T129 = T134 && T130;
  assign T130 = dramBank6_valid_received_1 || T131;
  assign T131 = dramBank6Port_rep_valid && T132;
  assign T132 = dramBank6Port_rep_tag == T133;
  assign T133 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T134 = ! T135;
  assign T135 = T136 == 5'h1/* 1*/;
  assign T136 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T137 = dramBank6_valid_received_0 & T138;
  assign T138 = T23[1'h0/* 0*/];
  assign T139 = T144 && T140;
  assign T140 = dramBank6_valid_received_0 || T141;
  assign T141 = dramBank6Port_rep_valid && T142;
  assign T142 = dramBank6Port_rep_tag == T143;
  assign T143 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T148 = ! dramBank6PortHadReadyRequest;
  assign T149 = T151 && T150;
  assign T150 = dramBank6PortHadReadyRequest || dramBank6Port_req_valid;
  assign T151 = ! AllOffloadsReady;
  assign T152 = dramBank6Port_req_ready || dramBank6_ready_received;
  assign T153 = T155 && T154;
  assign T154 = dramBank6_ready_received || dramBank6Port_req_ready;
  assign dramBank6Port_req_ready = mainOff_dramBank6_req_ready;
  assign T155 = ! AllOffloadsReady;
  assign T156 = T256 && T157;
  assign T157 = T252 || T158;
  assign T158 = T248 && T159;
  assign T159 = ! dramBank5Port_req_valid;
  assign dramBank5Port_req_valid = T160;
  assign T160 = T165 && T161;
  assign T161 = T164 && T162;
  assign T162 = T19 == T163;
  assign T163 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T164 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T165 = T247 && T166;
  assign T166 = ! T167;
  assign T167 = T178 | T168;
  assign T168 = dramBank5_valid_received_7 & T22;
  assign T169 = T175 && T170;
  assign T170 = dramBank5_valid_received_7 || T171;
  assign T171 = dramBank5Port_rep_valid && T172;
  assign T172 = dramBank5Port_rep_tag == T173;
  assign T173 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank5Port_rep_tag = mainOff_dramBank5_rep_tag;
  assign mainOff_dramBank5_rep_ready = dramBank5Port_rep_ready;
  assign dramBank5Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank5_req_valid = dramBank5Port_req_valid;
  assign mainOff_dramBank5_req_tag = dramBank5Port_req_tag;
  assign dramBank5Port_req_tag = T174;
  assign T174 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank5Port_rep_valid = mainOff_dramBank5_rep_valid;
  assign T175 = ! T176;
  assign T176 = T177 == 5'h7/* 7*/;
  assign T177 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T178 = T188 | T179;
  assign T179 = dramBank5_valid_received_6 & T73;
  assign T180 = T185 && T181;
  assign T181 = dramBank5_valid_received_6 || T182;
  assign T182 = dramBank5Port_rep_valid && T183;
  assign T183 = dramBank5Port_rep_tag == T184;
  assign T184 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T185 = ! T186;
  assign T186 = T187 == 5'h6/* 6*/;
  assign T187 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T188 = T198 | T189;
  assign T189 = dramBank5_valid_received_5 & T84;
  assign T190 = T195 && T191;
  assign T191 = dramBank5_valid_received_5 || T192;
  assign T192 = dramBank5Port_rep_valid && T193;
  assign T193 = dramBank5Port_rep_tag == T194;
  assign T194 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T195 = ! T196;
  assign T196 = T197 == 5'h5/* 5*/;
  assign T197 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T198 = T208 | T199;
  assign T199 = dramBank5_valid_received_4 & T95;
  assign T200 = T205 && T201;
  assign T201 = dramBank5_valid_received_4 || T202;
  assign T202 = dramBank5Port_rep_valid && T203;
  assign T203 = dramBank5Port_rep_tag == T204;
  assign T204 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T205 = ! T206;
  assign T206 = T207 == 5'h4/* 4*/;
  assign T207 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T208 = T218 | T209;
  assign T209 = dramBank5_valid_received_3 & T106;
  assign T210 = T215 && T211;
  assign T211 = dramBank5_valid_received_3 || T212;
  assign T212 = dramBank5Port_rep_valid && T213;
  assign T213 = dramBank5Port_rep_tag == T214;
  assign T214 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T215 = ! T216;
  assign T216 = T217 == 5'h3/* 3*/;
  assign T217 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T218 = T228 | T219;
  assign T219 = dramBank5_valid_received_2 & T117;
  assign T220 = T225 && T221;
  assign T221 = dramBank5_valid_received_2 || T222;
  assign T222 = dramBank5Port_rep_valid && T223;
  assign T223 = dramBank5Port_rep_tag == T224;
  assign T224 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T225 = ! T226;
  assign T226 = T227 == 5'h2/* 2*/;
  assign T227 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T228 = T238 | T229;
  assign T229 = dramBank5_valid_received_1 & T128;
  assign T230 = T235 && T231;
  assign T231 = dramBank5_valid_received_1 || T232;
  assign T232 = dramBank5Port_rep_valid && T233;
  assign T233 = dramBank5Port_rep_tag == T234;
  assign T234 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T235 = ! T236;
  assign T236 = T237 == 5'h1/* 1*/;
  assign T237 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T238 = dramBank5_valid_received_0 & T138;
  assign T239 = T244 && T240;
  assign T240 = dramBank5_valid_received_0 || T241;
  assign T241 = dramBank5Port_rep_valid && T242;
  assign T242 = dramBank5Port_rep_tag == T243;
  assign T243 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T244 = ! T245;
  assign T245 = T246 == 5'h0/* 0*/;
  assign T246 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T247 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T248 = ! dramBank5PortHadReadyRequest;
  assign T249 = T251 && T250;
  assign T250 = dramBank5PortHadReadyRequest || dramBank5Port_req_valid;
  assign T251 = ! AllOffloadsReady;
  assign T252 = dramBank5Port_req_ready || dramBank5_ready_received;
  assign T253 = T255 && T254;
  assign T254 = dramBank5_ready_received || dramBank5Port_req_ready;
  assign dramBank5Port_req_ready = mainOff_dramBank5_req_ready;
  assign T255 = ! AllOffloadsReady;
  assign T256 = T356 && T257;
  assign T257 = T352 || T258;
  assign T258 = T348 && T259;
  assign T259 = ! dramBank4Port_req_valid;
  assign dramBank4Port_req_valid = T260;
  assign T260 = T265 && T261;
  assign T261 = T264 && T262;
  assign T262 = T19 == T263;
  assign T263 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T264 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T265 = T347 && T266;
  assign T266 = ! T267;
  assign T267 = T278 | T268;
  assign T268 = dramBank4_valid_received_7 & T22;
  assign T269 = T275 && T270;
  assign T270 = dramBank4_valid_received_7 || T271;
  assign T271 = dramBank4Port_rep_valid && T272;
  assign T272 = dramBank4Port_rep_tag == T273;
  assign T273 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank4Port_rep_tag = mainOff_dramBank4_rep_tag;
  assign mainOff_dramBank4_rep_ready = dramBank4Port_rep_ready;
  assign dramBank4Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank4_req_valid = dramBank4Port_req_valid;
  assign mainOff_dramBank4_req_tag = dramBank4Port_req_tag;
  assign dramBank4Port_req_tag = T274;
  assign T274 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank4Port_rep_valid = mainOff_dramBank4_rep_valid;
  assign T275 = ! T276;
  assign T276 = T277 == 5'h7/* 7*/;
  assign T277 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T278 = T288 | T279;
  assign T279 = dramBank4_valid_received_6 & T73;
  assign T280 = T285 && T281;
  assign T281 = dramBank4_valid_received_6 || T282;
  assign T282 = dramBank4Port_rep_valid && T283;
  assign T283 = dramBank4Port_rep_tag == T284;
  assign T284 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T285 = ! T286;
  assign T286 = T287 == 5'h6/* 6*/;
  assign T287 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T288 = T298 | T289;
  assign T289 = dramBank4_valid_received_5 & T84;
  assign T290 = T295 && T291;
  assign T291 = dramBank4_valid_received_5 || T292;
  assign T292 = dramBank4Port_rep_valid && T293;
  assign T293 = dramBank4Port_rep_tag == T294;
  assign T294 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T295 = ! T296;
  assign T296 = T297 == 5'h5/* 5*/;
  assign T297 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T298 = T308 | T299;
  assign T299 = dramBank4_valid_received_4 & T95;
  assign T300 = T305 && T301;
  assign T301 = dramBank4_valid_received_4 || T302;
  assign T302 = dramBank4Port_rep_valid && T303;
  assign T303 = dramBank4Port_rep_tag == T304;
  assign T304 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T305 = ! T306;
  assign T306 = T307 == 5'h4/* 4*/;
  assign T307 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T308 = T318 | T309;
  assign T309 = dramBank4_valid_received_3 & T106;
  assign T310 = T315 && T311;
  assign T311 = dramBank4_valid_received_3 || T312;
  assign T312 = dramBank4Port_rep_valid && T313;
  assign T313 = dramBank4Port_rep_tag == T314;
  assign T314 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T315 = ! T316;
  assign T316 = T317 == 5'h3/* 3*/;
  assign T317 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T318 = T328 | T319;
  assign T319 = dramBank4_valid_received_2 & T117;
  assign T320 = T325 && T321;
  assign T321 = dramBank4_valid_received_2 || T322;
  assign T322 = dramBank4Port_rep_valid && T323;
  assign T323 = dramBank4Port_rep_tag == T324;
  assign T324 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T325 = ! T326;
  assign T326 = T327 == 5'h2/* 2*/;
  assign T327 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T328 = T338 | T329;
  assign T329 = dramBank4_valid_received_1 & T128;
  assign T330 = T335 && T331;
  assign T331 = dramBank4_valid_received_1 || T332;
  assign T332 = dramBank4Port_rep_valid && T333;
  assign T333 = dramBank4Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T335 = ! T336;
  assign T336 = T337 == 5'h1/* 1*/;
  assign T337 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T338 = dramBank4_valid_received_0 & T138;
  assign T339 = T344 && T340;
  assign T340 = dramBank4_valid_received_0 || T341;
  assign T341 = dramBank4Port_rep_valid && T342;
  assign T342 = dramBank4Port_rep_tag == T343;
  assign T343 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T344 = ! T345;
  assign T345 = T346 == 5'h0/* 0*/;
  assign T346 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T347 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T348 = ! dramBank4PortHadReadyRequest;
  assign T349 = T351 && T350;
  assign T350 = dramBank4PortHadReadyRequest || dramBank4Port_req_valid;
  assign T351 = ! AllOffloadsReady;
  assign T352 = dramBank4Port_req_ready || dramBank4_ready_received;
  assign T353 = T355 && T354;
  assign T354 = dramBank4_ready_received || dramBank4Port_req_ready;
  assign dramBank4Port_req_ready = mainOff_dramBank4_req_ready;
  assign T355 = ! AllOffloadsReady;
  assign T356 = T456 && T357;
  assign T357 = T452 || T358;
  assign T358 = T448 && T359;
  assign T359 = ! dramBank3Port_req_valid;
  assign dramBank3Port_req_valid = T360;
  assign T360 = T365 && T361;
  assign T361 = T364 && T362;
  assign T362 = T19 == T363;
  assign T363 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T364 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T365 = T447 && T366;
  assign T366 = ! T367;
  assign T367 = T378 | T368;
  assign T368 = dramBank3_valid_received_7 & T22;
  assign T369 = T375 && T370;
  assign T370 = dramBank3_valid_received_7 || T371;
  assign T371 = dramBank3Port_rep_valid && T372;
  assign T372 = dramBank3Port_rep_tag == T373;
  assign T373 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank3Port_rep_tag = mainOff_dramBank3_rep_tag;
  assign mainOff_dramBank3_rep_ready = dramBank3Port_rep_ready;
  assign dramBank3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank3_req_valid = dramBank3Port_req_valid;
  assign mainOff_dramBank3_req_tag = dramBank3Port_req_tag;
  assign dramBank3Port_req_tag = T374;
  assign T374 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank3Port_rep_valid = mainOff_dramBank3_rep_valid;
  assign T375 = ! T376;
  assign T376 = T377 == 5'h7/* 7*/;
  assign T377 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T378 = T388 | T379;
  assign T379 = dramBank3_valid_received_6 & T73;
  assign T380 = T385 && T381;
  assign T381 = dramBank3_valid_received_6 || T382;
  assign T382 = dramBank3Port_rep_valid && T383;
  assign T383 = dramBank3Port_rep_tag == T384;
  assign T384 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T385 = ! T386;
  assign T386 = T387 == 5'h6/* 6*/;
  assign T387 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T388 = T398 | T389;
  assign T389 = dramBank3_valid_received_5 & T84;
  assign T390 = T395 && T391;
  assign T391 = dramBank3_valid_received_5 || T392;
  assign T392 = dramBank3Port_rep_valid && T393;
  assign T393 = dramBank3Port_rep_tag == T394;
  assign T394 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T395 = ! T396;
  assign T396 = T397 == 5'h5/* 5*/;
  assign T397 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T398 = T408 | T399;
  assign T399 = dramBank3_valid_received_4 & T95;
  assign T400 = T405 && T401;
  assign T401 = dramBank3_valid_received_4 || T402;
  assign T402 = dramBank3Port_rep_valid && T403;
  assign T403 = dramBank3Port_rep_tag == T404;
  assign T404 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T405 = ! T406;
  assign T406 = T407 == 5'h4/* 4*/;
  assign T407 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T408 = T418 | T409;
  assign T409 = dramBank3_valid_received_3 & T106;
  assign T410 = T415 && T411;
  assign T411 = dramBank3_valid_received_3 || T412;
  assign T412 = dramBank3Port_rep_valid && T413;
  assign T413 = dramBank3Port_rep_tag == T414;
  assign T414 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T415 = ! T416;
  assign T416 = T417 == 5'h3/* 3*/;
  assign T417 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T418 = T428 | T419;
  assign T419 = dramBank3_valid_received_2 & T117;
  assign T420 = T425 && T421;
  assign T421 = dramBank3_valid_received_2 || T422;
  assign T422 = dramBank3Port_rep_valid && T423;
  assign T423 = dramBank3Port_rep_tag == T424;
  assign T424 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T425 = ! T426;
  assign T426 = T427 == 5'h2/* 2*/;
  assign T427 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T428 = T438 | T429;
  assign T429 = dramBank3_valid_received_1 & T128;
  assign T430 = T435 && T431;
  assign T431 = dramBank3_valid_received_1 || T432;
  assign T432 = dramBank3Port_rep_valid && T433;
  assign T433 = dramBank3Port_rep_tag == T434;
  assign T434 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T435 = ! T436;
  assign T436 = T437 == 5'h1/* 1*/;
  assign T437 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T438 = dramBank3_valid_received_0 & T138;
  assign T439 = T444 && T440;
  assign T440 = dramBank3_valid_received_0 || T441;
  assign T441 = dramBank3Port_rep_valid && T442;
  assign T442 = dramBank3Port_rep_tag == T443;
  assign T443 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T444 = ! T445;
  assign T445 = T446 == 5'h0/* 0*/;
  assign T446 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T447 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T448 = ! dramBank3PortHadReadyRequest;
  assign T449 = T451 && T450;
  assign T450 = dramBank3PortHadReadyRequest || dramBank3Port_req_valid;
  assign T451 = ! AllOffloadsReady;
  assign T452 = dramBank3Port_req_ready || dramBank3_ready_received;
  assign T453 = T455 && T454;
  assign T454 = dramBank3_ready_received || dramBank3Port_req_ready;
  assign dramBank3Port_req_ready = mainOff_dramBank3_req_ready;
  assign T455 = ! AllOffloadsReady;
  assign T456 = T556 && T457;
  assign T457 = T552 || T458;
  assign T458 = T548 && T459;
  assign T459 = ! dramBank2Port_req_valid;
  assign dramBank2Port_req_valid = T460;
  assign T460 = T465 && T461;
  assign T461 = T464 && T462;
  assign T462 = T19 == T463;
  assign T463 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T464 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T465 = T547 && T466;
  assign T466 = ! T467;
  assign T467 = T478 | T468;
  assign T468 = dramBank2_valid_received_7 & T22;
  assign T469 = T475 && T470;
  assign T470 = dramBank2_valid_received_7 || T471;
  assign T471 = dramBank2Port_rep_valid && T472;
  assign T472 = dramBank2Port_rep_tag == T473;
  assign T473 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank2Port_rep_tag = mainOff_dramBank2_rep_tag;
  assign mainOff_dramBank2_rep_ready = dramBank2Port_rep_ready;
  assign dramBank2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank2_req_valid = dramBank2Port_req_valid;
  assign mainOff_dramBank2_req_tag = dramBank2Port_req_tag;
  assign dramBank2Port_req_tag = T474;
  assign T474 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank2Port_rep_valid = mainOff_dramBank2_rep_valid;
  assign T475 = ! T476;
  assign T476 = T477 == 5'h7/* 7*/;
  assign T477 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T478 = T488 | T479;
  assign T479 = dramBank2_valid_received_6 & T73;
  assign T480 = T485 && T481;
  assign T481 = dramBank2_valid_received_6 || T482;
  assign T482 = dramBank2Port_rep_valid && T483;
  assign T483 = dramBank2Port_rep_tag == T484;
  assign T484 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T485 = ! T486;
  assign T486 = T487 == 5'h6/* 6*/;
  assign T487 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T488 = T498 | T489;
  assign T489 = dramBank2_valid_received_5 & T84;
  assign T490 = T495 && T491;
  assign T491 = dramBank2_valid_received_5 || T492;
  assign T492 = dramBank2Port_rep_valid && T493;
  assign T493 = dramBank2Port_rep_tag == T494;
  assign T494 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T495 = ! T496;
  assign T496 = T497 == 5'h5/* 5*/;
  assign T497 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T498 = T508 | T499;
  assign T499 = dramBank2_valid_received_4 & T95;
  assign T500 = T505 && T501;
  assign T501 = dramBank2_valid_received_4 || T502;
  assign T502 = dramBank2Port_rep_valid && T503;
  assign T503 = dramBank2Port_rep_tag == T504;
  assign T504 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T505 = ! T506;
  assign T506 = T507 == 5'h4/* 4*/;
  assign T507 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T508 = T518 | T509;
  assign T509 = dramBank2_valid_received_3 & T106;
  assign T510 = T515 && T511;
  assign T511 = dramBank2_valid_received_3 || T512;
  assign T512 = dramBank2Port_rep_valid && T513;
  assign T513 = dramBank2Port_rep_tag == T514;
  assign T514 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T515 = ! T516;
  assign T516 = T517 == 5'h3/* 3*/;
  assign T517 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T518 = T528 | T519;
  assign T519 = dramBank2_valid_received_2 & T117;
  assign T520 = T525 && T521;
  assign T521 = dramBank2_valid_received_2 || T522;
  assign T522 = dramBank2Port_rep_valid && T523;
  assign T523 = dramBank2Port_rep_tag == T524;
  assign T524 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T525 = ! T526;
  assign T526 = T527 == 5'h2/* 2*/;
  assign T527 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T528 = T538 | T529;
  assign T529 = dramBank2_valid_received_1 & T128;
  assign T530 = T535 && T531;
  assign T531 = dramBank2_valid_received_1 || T532;
  assign T532 = dramBank2Port_rep_valid && T533;
  assign T533 = dramBank2Port_rep_tag == T534;
  assign T534 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T535 = ! T536;
  assign T536 = T537 == 5'h1/* 1*/;
  assign T537 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T538 = dramBank2_valid_received_0 & T138;
  assign T539 = T544 && T540;
  assign T540 = dramBank2_valid_received_0 || T541;
  assign T541 = dramBank2Port_rep_valid && T542;
  assign T542 = dramBank2Port_rep_tag == T543;
  assign T543 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T544 = ! T545;
  assign T545 = T546 == 5'h0/* 0*/;
  assign T546 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T547 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T548 = ! dramBank2PortHadReadyRequest;
  assign T549 = T551 && T550;
  assign T550 = dramBank2PortHadReadyRequest || dramBank2Port_req_valid;
  assign T551 = ! AllOffloadsReady;
  assign T552 = dramBank2Port_req_ready || dramBank2_ready_received;
  assign T553 = T555 && T554;
  assign T554 = dramBank2_ready_received || dramBank2Port_req_ready;
  assign dramBank2Port_req_ready = mainOff_dramBank2_req_ready;
  assign T555 = ! AllOffloadsReady;
  assign T556 = T656 && T557;
  assign T557 = T652 || T558;
  assign T558 = T648 && T559;
  assign T559 = ! dramBank1Port_req_valid;
  assign dramBank1Port_req_valid = T560;
  assign T560 = T565 && T561;
  assign T561 = T564 && T562;
  assign T562 = T19 == T563;
  assign T563 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T564 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T565 = T647 && T566;
  assign T566 = ! T567;
  assign T567 = T578 | T568;
  assign T568 = dramBank1_valid_received_7 & T22;
  assign T569 = T575 && T570;
  assign T570 = dramBank1_valid_received_7 || T571;
  assign T571 = dramBank1Port_rep_valid && T572;
  assign T572 = dramBank1Port_rep_tag == T573;
  assign T573 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank1Port_rep_tag = mainOff_dramBank1_rep_tag;
  assign mainOff_dramBank1_rep_ready = dramBank1Port_rep_ready;
  assign dramBank1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank1_req_valid = dramBank1Port_req_valid;
  assign mainOff_dramBank1_req_tag = dramBank1Port_req_tag;
  assign dramBank1Port_req_tag = T574;
  assign T574 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank1Port_rep_valid = mainOff_dramBank1_rep_valid;
  assign T575 = ! T576;
  assign T576 = T577 == 5'h7/* 7*/;
  assign T577 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T578 = T588 | T579;
  assign T579 = dramBank1_valid_received_6 & T73;
  assign T580 = T585 && T581;
  assign T581 = dramBank1_valid_received_6 || T582;
  assign T582 = dramBank1Port_rep_valid && T583;
  assign T583 = dramBank1Port_rep_tag == T584;
  assign T584 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T585 = ! T586;
  assign T586 = T587 == 5'h6/* 6*/;
  assign T587 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T588 = T598 | T589;
  assign T589 = dramBank1_valid_received_5 & T84;
  assign T590 = T595 && T591;
  assign T591 = dramBank1_valid_received_5 || T592;
  assign T592 = dramBank1Port_rep_valid && T593;
  assign T593 = dramBank1Port_rep_tag == T594;
  assign T594 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T595 = ! T596;
  assign T596 = T597 == 5'h5/* 5*/;
  assign T597 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T598 = T608 | T599;
  assign T599 = dramBank1_valid_received_4 & T95;
  assign T600 = T605 && T601;
  assign T601 = dramBank1_valid_received_4 || T602;
  assign T602 = dramBank1Port_rep_valid && T603;
  assign T603 = dramBank1Port_rep_tag == T604;
  assign T604 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T605 = ! T606;
  assign T606 = T607 == 5'h4/* 4*/;
  assign T607 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T608 = T618 | T609;
  assign T609 = dramBank1_valid_received_3 & T106;
  assign T610 = T615 && T611;
  assign T611 = dramBank1_valid_received_3 || T612;
  assign T612 = dramBank1Port_rep_valid && T613;
  assign T613 = dramBank1Port_rep_tag == T614;
  assign T614 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T615 = ! T616;
  assign T616 = T617 == 5'h3/* 3*/;
  assign T617 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T618 = T628 | T619;
  assign T619 = dramBank1_valid_received_2 & T117;
  assign T620 = T625 && T621;
  assign T621 = dramBank1_valid_received_2 || T622;
  assign T622 = dramBank1Port_rep_valid && T623;
  assign T623 = dramBank1Port_rep_tag == T624;
  assign T624 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T625 = ! T626;
  assign T626 = T627 == 5'h2/* 2*/;
  assign T627 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T628 = T638 | T629;
  assign T629 = dramBank1_valid_received_1 & T128;
  assign T630 = T635 && T631;
  assign T631 = dramBank1_valid_received_1 || T632;
  assign T632 = dramBank1Port_rep_valid && T633;
  assign T633 = dramBank1Port_rep_tag == T634;
  assign T634 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T635 = ! T636;
  assign T636 = T637 == 5'h1/* 1*/;
  assign T637 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T638 = dramBank1_valid_received_0 & T138;
  assign T639 = T644 && T640;
  assign T640 = dramBank1_valid_received_0 || T641;
  assign T641 = dramBank1Port_rep_valid && T642;
  assign T642 = dramBank1Port_rep_tag == T643;
  assign T643 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T644 = ! T645;
  assign T645 = T646 == 5'h0/* 0*/;
  assign T646 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T647 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T648 = ! dramBank1PortHadReadyRequest;
  assign T649 = T651 && T650;
  assign T650 = dramBank1PortHadReadyRequest || dramBank1Port_req_valid;
  assign T651 = ! AllOffloadsReady;
  assign T652 = dramBank1Port_req_ready || dramBank1_ready_received;
  assign T653 = T655 && T654;
  assign T654 = dramBank1_ready_received || dramBank1Port_req_ready;
  assign dramBank1Port_req_ready = mainOff_dramBank1_req_ready;
  assign T655 = ! AllOffloadsReady;
  assign T656 = T751 || T657;
  assign T657 = T747 && T658;
  assign T658 = ! dramBank0Port_req_valid;
  assign dramBank0Port_req_valid = T659;
  assign T659 = T664 && T660;
  assign T660 = T663 && T661;
  assign T661 = T19 == T662;
  assign T662 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T663 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T664 = T746 && T665;
  assign T665 = ! T666;
  assign T666 = T677 | T667;
  assign T667 = dramBank0_valid_received_7 & T22;
  assign T668 = T674 && T669;
  assign T669 = dramBank0_valid_received_7 || T670;
  assign T670 = dramBank0Port_rep_valid && T671;
  assign T671 = dramBank0Port_rep_tag == T672;
  assign T672 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank0Port_rep_tag = mainOff_dramBank0_rep_tag;
  assign mainOff_dramBank0_rep_ready = dramBank0Port_rep_ready;
  assign dramBank0Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_dramBank0_req_valid = dramBank0Port_req_valid;
  assign mainOff_dramBank0_req_tag = dramBank0Port_req_tag;
  assign dramBank0Port_req_tag = T673;
  assign T673 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank0Port_rep_valid = mainOff_dramBank0_rep_valid;
  assign T674 = ! T675;
  assign T675 = T676 == 5'h7/* 7*/;
  assign T676 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T677 = T687 | T678;
  assign T678 = dramBank0_valid_received_6 & T73;
  assign T679 = T684 && T680;
  assign T680 = dramBank0_valid_received_6 || T681;
  assign T681 = dramBank0Port_rep_valid && T682;
  assign T682 = dramBank0Port_rep_tag == T683;
  assign T683 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T684 = ! T685;
  assign T685 = T686 == 5'h6/* 6*/;
  assign T686 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T687 = T697 | T688;
  assign T688 = dramBank0_valid_received_5 & T84;
  assign T689 = T694 && T690;
  assign T690 = dramBank0_valid_received_5 || T691;
  assign T691 = dramBank0Port_rep_valid && T692;
  assign T692 = dramBank0Port_rep_tag == T693;
  assign T693 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T694 = ! T695;
  assign T695 = T696 == 5'h5/* 5*/;
  assign T696 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T697 = T707 | T698;
  assign T698 = dramBank0_valid_received_4 & T95;
  assign T699 = T704 && T700;
  assign T700 = dramBank0_valid_received_4 || T701;
  assign T701 = dramBank0Port_rep_valid && T702;
  assign T702 = dramBank0Port_rep_tag == T703;
  assign T703 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T704 = ! T705;
  assign T705 = T706 == 5'h4/* 4*/;
  assign T706 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T707 = T717 | T708;
  assign T708 = dramBank0_valid_received_3 & T106;
  assign T709 = T714 && T710;
  assign T710 = dramBank0_valid_received_3 || T711;
  assign T711 = dramBank0Port_rep_valid && T712;
  assign T712 = dramBank0Port_rep_tag == T713;
  assign T713 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h3/* 3*/;
  assign T716 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T727 | T718;
  assign T718 = dramBank0_valid_received_2 & T117;
  assign T719 = T724 && T720;
  assign T720 = dramBank0_valid_received_2 || T721;
  assign T721 = dramBank0Port_rep_valid && T722;
  assign T722 = dramBank0Port_rep_tag == T723;
  assign T723 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T724 = ! T725;
  assign T725 = T726 == 5'h2/* 2*/;
  assign T726 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T727 = T737 | T728;
  assign T728 = dramBank0_valid_received_1 & T128;
  assign T729 = T734 && T730;
  assign T730 = dramBank0_valid_received_1 || T731;
  assign T731 = dramBank0Port_rep_valid && T732;
  assign T732 = dramBank0Port_rep_tag == T733;
  assign T733 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T734 = ! T735;
  assign T735 = T736 == 5'h1/* 1*/;
  assign T736 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T737 = dramBank0_valid_received_0 & T138;
  assign T738 = T743 && T739;
  assign T739 = dramBank0_valid_received_0 || T740;
  assign T740 = dramBank0Port_rep_valid && T741;
  assign T741 = dramBank0Port_rep_tag == T742;
  assign T742 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h0/* 0*/;
  assign T745 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T747 = ! dramBank0PortHadReadyRequest;
  assign T748 = T750 && T749;
  assign T749 = dramBank0PortHadReadyRequest || dramBank0Port_req_valid;
  assign T750 = ! AllOffloadsReady;
  assign T751 = dramBank0Port_req_ready || dramBank0_ready_received;
  assign T752 = T754 && T753;
  assign T753 = dramBank0_ready_received || dramBank0Port_req_ready;
  assign dramBank0Port_req_ready = mainOff_dramBank0_req_ready;
  assign T754 = ! AllOffloadsReady;
  assign T755 = subStateTh_6 == 1'h0/* 0*/;
  assign T756 = T760 ? 1'h1/* 1*/ : T757;
  assign T757 = T758 ? 1'h0/* 0*/ : subStateTh_6;
  assign T758 = T759 == vThreadEncoder_io_chosen;
  assign T759 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T760 = T2286 && T761;
  assign T761 = State_6 != 8'hff/* 255*/;
  assign T762 = T2204 || T763;
  assign T763 = T765 && T764;
  assign T764 = T6[3'h6/* 6*/];
  assign T765 = T2203 && T766;
  assign T766 = T768 == T767;
  assign T767 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T768 = T771 | T769;
  assign T769 = State_7 & T770;
  assign T770 = {4'h8/* 8*/{T5}};
  assign T771 = T774 | T772;
  assign T772 = State_6 & T773;
  assign T773 = {4'h8/* 8*/{T764}};
  assign T774 = T1774 | T775;
  assign T775 = State_5 & T776;
  assign T776 = {4'h8/* 8*/{T777}};
  assign T777 = T6[3'h5/* 5*/];
  assign T778 = T780 || T779;
  assign T779 = T765 && T777;
  assign T780 = T786 || T781;
  assign T781 = T782 && T777;
  assign T782 = T785 && T783;
  assign T783 = T768 == T784;
  assign T784 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T785 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T786 = T792 || T787;
  assign T787 = T788 && T777;
  assign T788 = T791 && T789;
  assign T789 = T768 == T790;
  assign T790 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T791 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T792 = T798 || T793;
  assign T793 = T794 && T777;
  assign T794 = T797 && T795;
  assign T795 = T768 == T796;
  assign T796 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T797 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T798 = T804 || T799;
  assign T799 = T800 && T777;
  assign T800 = T803 && T801;
  assign T801 = T768 == T802;
  assign T802 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T803 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T804 = T810 || T805;
  assign T805 = T806 && T777;
  assign T806 = T809 && T807;
  assign T807 = T768 == T808;
  assign T808 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T809 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T810 = T816 || T811;
  assign T811 = T812 && T777;
  assign T812 = T815 && T813;
  assign T813 = T768 == T814;
  assign T814 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T815 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T816 = T822 || T817;
  assign T817 = T818 && T777;
  assign T818 = T821 && T819;
  assign T819 = T768 == T820;
  assign T820 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T821 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T822 = T828 || T823;
  assign T823 = T824 && T777;
  assign T824 = T827 && T825;
  assign T825 = T768 == T826;
  assign T826 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T827 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T828 = T924 || T829;
  assign T829 = T830 && T777;
  assign T830 = T892 && T831;
  assign T831 = ! T832;
  assign T832 = b == T833;
  assign T833 = {16'h0/* 0*/, 32'h7/* 7*/};
  assign b = T834 & 48'h7fff/* 32767*/;
  assign T834 = {16'h0/* 0*/, T835};
  assign T835 = T836 >> 33'hc/* 12*/;
  assign T836 = T846 | T837;
  assign T837 = inputReg_7_addr & T838;
  assign T838 = {6'h20/* 32*/{T5}};
  assign T839 = T843 && T840;
  assign T840 = T841[3'h7/* 7*/];
  assign T841 = T842[3'h7/* 7*/:1'h0/* 0*/];
  assign T842 = 8'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T843 = T844 && io_in_valid;
  assign T844 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T845 = T839 ? io_in_bits_addr : inputReg_7_addr;
  assign T846 = T852 | T847;
  assign T847 = inputReg_6_addr & T848;
  assign T848 = {6'h20/* 32*/{T764}};
  assign T849 = T843 && T850;
  assign T850 = T841[3'h6/* 6*/];
  assign T851 = T849 ? io_in_bits_addr : inputReg_6_addr;
  assign T852 = T858 | T853;
  assign T853 = inputReg_5_addr & T854;
  assign T854 = {6'h20/* 32*/{T777}};
  assign T855 = T843 && T856;
  assign T856 = T841[3'h5/* 5*/];
  assign T857 = T855 ? io_in_bits_addr : inputReg_5_addr;
  assign T858 = T865 | T859;
  assign T859 = inputReg_4_addr & T860;
  assign T860 = {6'h20/* 32*/{T861}};
  assign T861 = T6[3'h4/* 4*/];
  assign T862 = T843 && T863;
  assign T863 = T841[3'h4/* 4*/];
  assign T864 = T862 ? io_in_bits_addr : inputReg_4_addr;
  assign T865 = T872 | T866;
  assign T866 = inputReg_3_addr & T867;
  assign T867 = {6'h20/* 32*/{T868}};
  assign T868 = T6[2'h3/* 3*/];
  assign T869 = T843 && T870;
  assign T870 = T841[2'h3/* 3*/];
  assign T871 = T869 ? io_in_bits_addr : inputReg_3_addr;
  assign T872 = T879 | T873;
  assign T873 = inputReg_2_addr & T874;
  assign T874 = {6'h20/* 32*/{T875}};
  assign T875 = T6[2'h2/* 2*/];
  assign T876 = T843 && T877;
  assign T877 = T841[2'h2/* 2*/];
  assign T878 = T876 ? io_in_bits_addr : inputReg_2_addr;
  assign T879 = T886 | T880;
  assign T880 = inputReg_1_addr & T881;
  assign T881 = {6'h20/* 32*/{T882}};
  assign T882 = T6[1'h1/* 1*/];
  assign T883 = T843 && T884;
  assign T884 = T841[1'h1/* 1*/];
  assign T885 = T883 ? io_in_bits_addr : inputReg_1_addr;
  assign T886 = inputReg_0_addr & T887;
  assign T887 = {6'h20/* 32*/{T888}};
  assign T888 = T6[1'h0/* 0*/];
  assign T889 = T843 && T890;
  assign T890 = T841[1'h0/* 0*/];
  assign T891 = T889 ? io_in_bits_addr : inputReg_0_addr;
  assign T892 = T896 && T893;
  assign T893 = ! T894;
  assign T894 = b == T895;
  assign T895 = {16'h0/* 0*/, 32'h6/* 6*/};
  assign T896 = T900 && T897;
  assign T897 = ! T898;
  assign T898 = b == T899;
  assign T899 = {16'h0/* 0*/, 32'h5/* 5*/};
  assign T900 = T904 && T901;
  assign T901 = ! T902;
  assign T902 = b == T903;
  assign T903 = {16'h0/* 0*/, 32'h4/* 4*/};
  assign T904 = T908 && T905;
  assign T905 = ! T906;
  assign T906 = b == T907;
  assign T907 = {16'h0/* 0*/, 32'h3/* 3*/};
  assign T908 = T912 && T909;
  assign T909 = ! T910;
  assign T910 = b == T911;
  assign T911 = {16'h0/* 0*/, 32'h2/* 2*/};
  assign T912 = T916 && T913;
  assign T913 = ! T914;
  assign T914 = b == T915;
  assign T915 = {16'h0/* 0*/, 32'h1/* 1*/};
  assign T916 = T920 && T917;
  assign T917 = ! T918;
  assign T918 = b == T919;
  assign T919 = {16'h0/* 0*/, 32'h0/* 0*/};
  assign T920 = T923 && T921;
  assign T921 = T768 == T922;
  assign T922 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T923 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T924 = T995 || T925;
  assign T925 = T926 && T777;
  assign T926 = T994 && T927;
  assign T927 = ! T928;
  assign T928 = T931 == r;
  assign r = T929 & 60'h7ffffff/* 134217727*/;
  assign T929 = {28'h0/* 0*/, T930};
  assign T930 = T836 >> 34'hf/* 15*/;
  assign T931 = {28'h0/* 0*/, T932};
  assign T932 = T940 | T933;
  assign T933 = rb7RowAddr_7 & T934;
  assign T934 = {6'h20/* 32*/{T5}};
  assign T935 = T839 || T936;
  assign T936 = T926 && T5;
  assign T937 = T936 ? r : T938;
  assign T938 = {28'h0/* 0*/, T939};
  assign T939 = T839 ? 32'h0/* 0*/ : rb7RowAddr_7;
  assign T940 = T948 | T941;
  assign T941 = rb7RowAddr_6 & T942;
  assign T942 = {6'h20/* 32*/{T764}};
  assign T943 = T849 || T944;
  assign T944 = T926 && T764;
  assign T945 = T944 ? r : T946;
  assign T946 = {28'h0/* 0*/, T947};
  assign T947 = T849 ? 32'h0/* 0*/ : rb7RowAddr_6;
  assign T948 = T955 | T949;
  assign T949 = rb7RowAddr_5 & T950;
  assign T950 = {6'h20/* 32*/{T777}};
  assign T951 = T855 || T925;
  assign T952 = T925 ? r : T953;
  assign T953 = {28'h0/* 0*/, T954};
  assign T954 = T855 ? 32'h0/* 0*/ : rb7RowAddr_5;
  assign T955 = T963 | T956;
  assign T956 = rb7RowAddr_4 & T957;
  assign T957 = {6'h20/* 32*/{T861}};
  assign T958 = T862 || T959;
  assign T959 = T926 && T861;
  assign T960 = T959 ? r : T961;
  assign T961 = {28'h0/* 0*/, T962};
  assign T962 = T862 ? 32'h0/* 0*/ : rb7RowAddr_4;
  assign T963 = T971 | T964;
  assign T964 = rb7RowAddr_3 & T965;
  assign T965 = {6'h20/* 32*/{T868}};
  assign T966 = T869 || T967;
  assign T967 = T926 && T868;
  assign T968 = T967 ? r : T969;
  assign T969 = {28'h0/* 0*/, T970};
  assign T970 = T869 ? 32'h0/* 0*/ : rb7RowAddr_3;
  assign T971 = T979 | T972;
  assign T972 = rb7RowAddr_2 & T973;
  assign T973 = {6'h20/* 32*/{T875}};
  assign T974 = T876 || T975;
  assign T975 = T926 && T875;
  assign T976 = T975 ? r : T977;
  assign T977 = {28'h0/* 0*/, T978};
  assign T978 = T876 ? 32'h0/* 0*/ : rb7RowAddr_2;
  assign T979 = T987 | T980;
  assign T980 = rb7RowAddr_1 & T981;
  assign T981 = {6'h20/* 32*/{T882}};
  assign T982 = T883 || T983;
  assign T983 = T926 && T882;
  assign T984 = T983 ? r : T985;
  assign T985 = {28'h0/* 0*/, T986};
  assign T986 = T883 ? 32'h0/* 0*/ : rb7RowAddr_1;
  assign T987 = rb7RowAddr_0 & T988;
  assign T988 = {6'h20/* 32*/{T888}};
  assign T989 = T889 || T990;
  assign T990 = T926 && T888;
  assign T991 = T990 ? r : T992;
  assign T992 = {28'h0/* 0*/, T993};
  assign T993 = T889 ? 32'h0/* 0*/ : rb7RowAddr_0;
  assign T994 = T892 && T832;
  assign T995 = T998 || T996;
  assign T996 = T997 && T777;
  assign T997 = T994 && T928;
  assign T998 = T1067 || T999;
  assign T999 = T1000 && T777;
  assign T1000 = T1066 && T1001;
  assign T1001 = ! T1002;
  assign T1002 = T1003 == r;
  assign T1003 = {28'h0/* 0*/, T1004};
  assign T1004 = T1012 | T1005;
  assign T1005 = rb6RowAddr_7 & T1006;
  assign T1006 = {6'h20/* 32*/{T5}};
  assign T1007 = T839 || T1008;
  assign T1008 = T1000 && T5;
  assign T1009 = T1008 ? r : T1010;
  assign T1010 = {28'h0/* 0*/, T1011};
  assign T1011 = T839 ? 32'h0/* 0*/ : rb6RowAddr_7;
  assign T1012 = T1020 | T1013;
  assign T1013 = rb6RowAddr_6 & T1014;
  assign T1014 = {6'h20/* 32*/{T764}};
  assign T1015 = T849 || T1016;
  assign T1016 = T1000 && T764;
  assign T1017 = T1016 ? r : T1018;
  assign T1018 = {28'h0/* 0*/, T1019};
  assign T1019 = T849 ? 32'h0/* 0*/ : rb6RowAddr_6;
  assign T1020 = T1027 | T1021;
  assign T1021 = rb6RowAddr_5 & T1022;
  assign T1022 = {6'h20/* 32*/{T777}};
  assign T1023 = T855 || T999;
  assign T1024 = T999 ? r : T1025;
  assign T1025 = {28'h0/* 0*/, T1026};
  assign T1026 = T855 ? 32'h0/* 0*/ : rb6RowAddr_5;
  assign T1027 = T1035 | T1028;
  assign T1028 = rb6RowAddr_4 & T1029;
  assign T1029 = {6'h20/* 32*/{T861}};
  assign T1030 = T862 || T1031;
  assign T1031 = T1000 && T861;
  assign T1032 = T1031 ? r : T1033;
  assign T1033 = {28'h0/* 0*/, T1034};
  assign T1034 = T862 ? 32'h0/* 0*/ : rb6RowAddr_4;
  assign T1035 = T1043 | T1036;
  assign T1036 = rb6RowAddr_3 & T1037;
  assign T1037 = {6'h20/* 32*/{T868}};
  assign T1038 = T869 || T1039;
  assign T1039 = T1000 && T868;
  assign T1040 = T1039 ? r : T1041;
  assign T1041 = {28'h0/* 0*/, T1042};
  assign T1042 = T869 ? 32'h0/* 0*/ : rb6RowAddr_3;
  assign T1043 = T1051 | T1044;
  assign T1044 = rb6RowAddr_2 & T1045;
  assign T1045 = {6'h20/* 32*/{T875}};
  assign T1046 = T876 || T1047;
  assign T1047 = T1000 && T875;
  assign T1048 = T1047 ? r : T1049;
  assign T1049 = {28'h0/* 0*/, T1050};
  assign T1050 = T876 ? 32'h0/* 0*/ : rb6RowAddr_2;
  assign T1051 = T1059 | T1052;
  assign T1052 = rb6RowAddr_1 & T1053;
  assign T1053 = {6'h20/* 32*/{T882}};
  assign T1054 = T883 || T1055;
  assign T1055 = T1000 && T882;
  assign T1056 = T1055 ? r : T1057;
  assign T1057 = {28'h0/* 0*/, T1058};
  assign T1058 = T883 ? 32'h0/* 0*/ : rb6RowAddr_1;
  assign T1059 = rb6RowAddr_0 & T1060;
  assign T1060 = {6'h20/* 32*/{T888}};
  assign T1061 = T889 || T1062;
  assign T1062 = T1000 && T888;
  assign T1063 = T1062 ? r : T1064;
  assign T1064 = {28'h0/* 0*/, T1065};
  assign T1065 = T889 ? 32'h0/* 0*/ : rb6RowAddr_0;
  assign T1066 = T896 && T894;
  assign T1067 = T1070 || T1068;
  assign T1068 = T1069 && T777;
  assign T1069 = T1066 && T1002;
  assign T1070 = T1139 || T1071;
  assign T1071 = T1072 && T777;
  assign T1072 = T1138 && T1073;
  assign T1073 = ! T1074;
  assign T1074 = T1075 == r;
  assign T1075 = {28'h0/* 0*/, T1076};
  assign T1076 = T1084 | T1077;
  assign T1077 = rb5RowAddr_7 & T1078;
  assign T1078 = {6'h20/* 32*/{T5}};
  assign T1079 = T839 || T1080;
  assign T1080 = T1072 && T5;
  assign T1081 = T1080 ? r : T1082;
  assign T1082 = {28'h0/* 0*/, T1083};
  assign T1083 = T839 ? 32'h0/* 0*/ : rb5RowAddr_7;
  assign T1084 = T1092 | T1085;
  assign T1085 = rb5RowAddr_6 & T1086;
  assign T1086 = {6'h20/* 32*/{T764}};
  assign T1087 = T849 || T1088;
  assign T1088 = T1072 && T764;
  assign T1089 = T1088 ? r : T1090;
  assign T1090 = {28'h0/* 0*/, T1091};
  assign T1091 = T849 ? 32'h0/* 0*/ : rb5RowAddr_6;
  assign T1092 = T1099 | T1093;
  assign T1093 = rb5RowAddr_5 & T1094;
  assign T1094 = {6'h20/* 32*/{T777}};
  assign T1095 = T855 || T1071;
  assign T1096 = T1071 ? r : T1097;
  assign T1097 = {28'h0/* 0*/, T1098};
  assign T1098 = T855 ? 32'h0/* 0*/ : rb5RowAddr_5;
  assign T1099 = T1107 | T1100;
  assign T1100 = rb5RowAddr_4 & T1101;
  assign T1101 = {6'h20/* 32*/{T861}};
  assign T1102 = T862 || T1103;
  assign T1103 = T1072 && T861;
  assign T1104 = T1103 ? r : T1105;
  assign T1105 = {28'h0/* 0*/, T1106};
  assign T1106 = T862 ? 32'h0/* 0*/ : rb5RowAddr_4;
  assign T1107 = T1115 | T1108;
  assign T1108 = rb5RowAddr_3 & T1109;
  assign T1109 = {6'h20/* 32*/{T868}};
  assign T1110 = T869 || T1111;
  assign T1111 = T1072 && T868;
  assign T1112 = T1111 ? r : T1113;
  assign T1113 = {28'h0/* 0*/, T1114};
  assign T1114 = T869 ? 32'h0/* 0*/ : rb5RowAddr_3;
  assign T1115 = T1123 | T1116;
  assign T1116 = rb5RowAddr_2 & T1117;
  assign T1117 = {6'h20/* 32*/{T875}};
  assign T1118 = T876 || T1119;
  assign T1119 = T1072 && T875;
  assign T1120 = T1119 ? r : T1121;
  assign T1121 = {28'h0/* 0*/, T1122};
  assign T1122 = T876 ? 32'h0/* 0*/ : rb5RowAddr_2;
  assign T1123 = T1131 | T1124;
  assign T1124 = rb5RowAddr_1 & T1125;
  assign T1125 = {6'h20/* 32*/{T882}};
  assign T1126 = T883 || T1127;
  assign T1127 = T1072 && T882;
  assign T1128 = T1127 ? r : T1129;
  assign T1129 = {28'h0/* 0*/, T1130};
  assign T1130 = T883 ? 32'h0/* 0*/ : rb5RowAddr_1;
  assign T1131 = rb5RowAddr_0 & T1132;
  assign T1132 = {6'h20/* 32*/{T888}};
  assign T1133 = T889 || T1134;
  assign T1134 = T1072 && T888;
  assign T1135 = T1134 ? r : T1136;
  assign T1136 = {28'h0/* 0*/, T1137};
  assign T1137 = T889 ? 32'h0/* 0*/ : rb5RowAddr_0;
  assign T1138 = T900 && T898;
  assign T1139 = T1142 || T1140;
  assign T1140 = T1141 && T777;
  assign T1141 = T1138 && T1074;
  assign T1142 = T1211 || T1143;
  assign T1143 = T1144 && T777;
  assign T1144 = T1210 && T1145;
  assign T1145 = ! T1146;
  assign T1146 = T1147 == r;
  assign T1147 = {28'h0/* 0*/, T1148};
  assign T1148 = T1156 | T1149;
  assign T1149 = rb4RowAddr_7 & T1150;
  assign T1150 = {6'h20/* 32*/{T5}};
  assign T1151 = T839 || T1152;
  assign T1152 = T1144 && T5;
  assign T1153 = T1152 ? r : T1154;
  assign T1154 = {28'h0/* 0*/, T1155};
  assign T1155 = T839 ? 32'h0/* 0*/ : rb4RowAddr_7;
  assign T1156 = T1164 | T1157;
  assign T1157 = rb4RowAddr_6 & T1158;
  assign T1158 = {6'h20/* 32*/{T764}};
  assign T1159 = T849 || T1160;
  assign T1160 = T1144 && T764;
  assign T1161 = T1160 ? r : T1162;
  assign T1162 = {28'h0/* 0*/, T1163};
  assign T1163 = T849 ? 32'h0/* 0*/ : rb4RowAddr_6;
  assign T1164 = T1171 | T1165;
  assign T1165 = rb4RowAddr_5 & T1166;
  assign T1166 = {6'h20/* 32*/{T777}};
  assign T1167 = T855 || T1143;
  assign T1168 = T1143 ? r : T1169;
  assign T1169 = {28'h0/* 0*/, T1170};
  assign T1170 = T855 ? 32'h0/* 0*/ : rb4RowAddr_5;
  assign T1171 = T1179 | T1172;
  assign T1172 = rb4RowAddr_4 & T1173;
  assign T1173 = {6'h20/* 32*/{T861}};
  assign T1174 = T862 || T1175;
  assign T1175 = T1144 && T861;
  assign T1176 = T1175 ? r : T1177;
  assign T1177 = {28'h0/* 0*/, T1178};
  assign T1178 = T862 ? 32'h0/* 0*/ : rb4RowAddr_4;
  assign T1179 = T1187 | T1180;
  assign T1180 = rb4RowAddr_3 & T1181;
  assign T1181 = {6'h20/* 32*/{T868}};
  assign T1182 = T869 || T1183;
  assign T1183 = T1144 && T868;
  assign T1184 = T1183 ? r : T1185;
  assign T1185 = {28'h0/* 0*/, T1186};
  assign T1186 = T869 ? 32'h0/* 0*/ : rb4RowAddr_3;
  assign T1187 = T1195 | T1188;
  assign T1188 = rb4RowAddr_2 & T1189;
  assign T1189 = {6'h20/* 32*/{T875}};
  assign T1190 = T876 || T1191;
  assign T1191 = T1144 && T875;
  assign T1192 = T1191 ? r : T1193;
  assign T1193 = {28'h0/* 0*/, T1194};
  assign T1194 = T876 ? 32'h0/* 0*/ : rb4RowAddr_2;
  assign T1195 = T1203 | T1196;
  assign T1196 = rb4RowAddr_1 & T1197;
  assign T1197 = {6'h20/* 32*/{T882}};
  assign T1198 = T883 || T1199;
  assign T1199 = T1144 && T882;
  assign T1200 = T1199 ? r : T1201;
  assign T1201 = {28'h0/* 0*/, T1202};
  assign T1202 = T883 ? 32'h0/* 0*/ : rb4RowAddr_1;
  assign T1203 = rb4RowAddr_0 & T1204;
  assign T1204 = {6'h20/* 32*/{T888}};
  assign T1205 = T889 || T1206;
  assign T1206 = T1144 && T888;
  assign T1207 = T1206 ? r : T1208;
  assign T1208 = {28'h0/* 0*/, T1209};
  assign T1209 = T889 ? 32'h0/* 0*/ : rb4RowAddr_0;
  assign T1210 = T904 && T902;
  assign T1211 = T1214 || T1212;
  assign T1212 = T1213 && T777;
  assign T1213 = T1210 && T1146;
  assign T1214 = T1283 || T1215;
  assign T1215 = T1216 && T777;
  assign T1216 = T1282 && T1217;
  assign T1217 = ! T1218;
  assign T1218 = T1219 == r;
  assign T1219 = {28'h0/* 0*/, T1220};
  assign T1220 = T1228 | T1221;
  assign T1221 = rb3RowAddr_7 & T1222;
  assign T1222 = {6'h20/* 32*/{T5}};
  assign T1223 = T839 || T1224;
  assign T1224 = T1216 && T5;
  assign T1225 = T1224 ? r : T1226;
  assign T1226 = {28'h0/* 0*/, T1227};
  assign T1227 = T839 ? 32'h0/* 0*/ : rb3RowAddr_7;
  assign T1228 = T1236 | T1229;
  assign T1229 = rb3RowAddr_6 & T1230;
  assign T1230 = {6'h20/* 32*/{T764}};
  assign T1231 = T849 || T1232;
  assign T1232 = T1216 && T764;
  assign T1233 = T1232 ? r : T1234;
  assign T1234 = {28'h0/* 0*/, T1235};
  assign T1235 = T849 ? 32'h0/* 0*/ : rb3RowAddr_6;
  assign T1236 = T1243 | T1237;
  assign T1237 = rb3RowAddr_5 & T1238;
  assign T1238 = {6'h20/* 32*/{T777}};
  assign T1239 = T855 || T1215;
  assign T1240 = T1215 ? r : T1241;
  assign T1241 = {28'h0/* 0*/, T1242};
  assign T1242 = T855 ? 32'h0/* 0*/ : rb3RowAddr_5;
  assign T1243 = T1251 | T1244;
  assign T1244 = rb3RowAddr_4 & T1245;
  assign T1245 = {6'h20/* 32*/{T861}};
  assign T1246 = T862 || T1247;
  assign T1247 = T1216 && T861;
  assign T1248 = T1247 ? r : T1249;
  assign T1249 = {28'h0/* 0*/, T1250};
  assign T1250 = T862 ? 32'h0/* 0*/ : rb3RowAddr_4;
  assign T1251 = T1259 | T1252;
  assign T1252 = rb3RowAddr_3 & T1253;
  assign T1253 = {6'h20/* 32*/{T868}};
  assign T1254 = T869 || T1255;
  assign T1255 = T1216 && T868;
  assign T1256 = T1255 ? r : T1257;
  assign T1257 = {28'h0/* 0*/, T1258};
  assign T1258 = T869 ? 32'h0/* 0*/ : rb3RowAddr_3;
  assign T1259 = T1267 | T1260;
  assign T1260 = rb3RowAddr_2 & T1261;
  assign T1261 = {6'h20/* 32*/{T875}};
  assign T1262 = T876 || T1263;
  assign T1263 = T1216 && T875;
  assign T1264 = T1263 ? r : T1265;
  assign T1265 = {28'h0/* 0*/, T1266};
  assign T1266 = T876 ? 32'h0/* 0*/ : rb3RowAddr_2;
  assign T1267 = T1275 | T1268;
  assign T1268 = rb3RowAddr_1 & T1269;
  assign T1269 = {6'h20/* 32*/{T882}};
  assign T1270 = T883 || T1271;
  assign T1271 = T1216 && T882;
  assign T1272 = T1271 ? r : T1273;
  assign T1273 = {28'h0/* 0*/, T1274};
  assign T1274 = T883 ? 32'h0/* 0*/ : rb3RowAddr_1;
  assign T1275 = rb3RowAddr_0 & T1276;
  assign T1276 = {6'h20/* 32*/{T888}};
  assign T1277 = T889 || T1278;
  assign T1278 = T1216 && T888;
  assign T1279 = T1278 ? r : T1280;
  assign T1280 = {28'h0/* 0*/, T1281};
  assign T1281 = T889 ? 32'h0/* 0*/ : rb3RowAddr_0;
  assign T1282 = T908 && T906;
  assign T1283 = T1286 || T1284;
  assign T1284 = T1285 && T777;
  assign T1285 = T1282 && T1218;
  assign T1286 = T1355 || T1287;
  assign T1287 = T1288 && T777;
  assign T1288 = T1354 && T1289;
  assign T1289 = ! T1290;
  assign T1290 = T1291 == r;
  assign T1291 = {28'h0/* 0*/, T1292};
  assign T1292 = T1300 | T1293;
  assign T1293 = rb2RowAddr_7 & T1294;
  assign T1294 = {6'h20/* 32*/{T5}};
  assign T1295 = T839 || T1296;
  assign T1296 = T1288 && T5;
  assign T1297 = T1296 ? r : T1298;
  assign T1298 = {28'h0/* 0*/, T1299};
  assign T1299 = T839 ? 32'h0/* 0*/ : rb2RowAddr_7;
  assign T1300 = T1308 | T1301;
  assign T1301 = rb2RowAddr_6 & T1302;
  assign T1302 = {6'h20/* 32*/{T764}};
  assign T1303 = T849 || T1304;
  assign T1304 = T1288 && T764;
  assign T1305 = T1304 ? r : T1306;
  assign T1306 = {28'h0/* 0*/, T1307};
  assign T1307 = T849 ? 32'h0/* 0*/ : rb2RowAddr_6;
  assign T1308 = T1315 | T1309;
  assign T1309 = rb2RowAddr_5 & T1310;
  assign T1310 = {6'h20/* 32*/{T777}};
  assign T1311 = T855 || T1287;
  assign T1312 = T1287 ? r : T1313;
  assign T1313 = {28'h0/* 0*/, T1314};
  assign T1314 = T855 ? 32'h0/* 0*/ : rb2RowAddr_5;
  assign T1315 = T1323 | T1316;
  assign T1316 = rb2RowAddr_4 & T1317;
  assign T1317 = {6'h20/* 32*/{T861}};
  assign T1318 = T862 || T1319;
  assign T1319 = T1288 && T861;
  assign T1320 = T1319 ? r : T1321;
  assign T1321 = {28'h0/* 0*/, T1322};
  assign T1322 = T862 ? 32'h0/* 0*/ : rb2RowAddr_4;
  assign T1323 = T1331 | T1324;
  assign T1324 = rb2RowAddr_3 & T1325;
  assign T1325 = {6'h20/* 32*/{T868}};
  assign T1326 = T869 || T1327;
  assign T1327 = T1288 && T868;
  assign T1328 = T1327 ? r : T1329;
  assign T1329 = {28'h0/* 0*/, T1330};
  assign T1330 = T869 ? 32'h0/* 0*/ : rb2RowAddr_3;
  assign T1331 = T1339 | T1332;
  assign T1332 = rb2RowAddr_2 & T1333;
  assign T1333 = {6'h20/* 32*/{T875}};
  assign T1334 = T876 || T1335;
  assign T1335 = T1288 && T875;
  assign T1336 = T1335 ? r : T1337;
  assign T1337 = {28'h0/* 0*/, T1338};
  assign T1338 = T876 ? 32'h0/* 0*/ : rb2RowAddr_2;
  assign T1339 = T1347 | T1340;
  assign T1340 = rb2RowAddr_1 & T1341;
  assign T1341 = {6'h20/* 32*/{T882}};
  assign T1342 = T883 || T1343;
  assign T1343 = T1288 && T882;
  assign T1344 = T1343 ? r : T1345;
  assign T1345 = {28'h0/* 0*/, T1346};
  assign T1346 = T883 ? 32'h0/* 0*/ : rb2RowAddr_1;
  assign T1347 = rb2RowAddr_0 & T1348;
  assign T1348 = {6'h20/* 32*/{T888}};
  assign T1349 = T889 || T1350;
  assign T1350 = T1288 && T888;
  assign T1351 = T1350 ? r : T1352;
  assign T1352 = {28'h0/* 0*/, T1353};
  assign T1353 = T889 ? 32'h0/* 0*/ : rb2RowAddr_0;
  assign T1354 = T912 && T910;
  assign T1355 = T1358 || T1356;
  assign T1356 = T1357 && T777;
  assign T1357 = T1354 && T1290;
  assign T1358 = T1427 || T1359;
  assign T1359 = T1360 && T777;
  assign T1360 = T1426 && T1361;
  assign T1361 = ! T1362;
  assign T1362 = T1363 == r;
  assign T1363 = {28'h0/* 0*/, T1364};
  assign T1364 = T1372 | T1365;
  assign T1365 = rb1RowAddr_7 & T1366;
  assign T1366 = {6'h20/* 32*/{T5}};
  assign T1367 = T839 || T1368;
  assign T1368 = T1360 && T5;
  assign T1369 = T1368 ? r : T1370;
  assign T1370 = {28'h0/* 0*/, T1371};
  assign T1371 = T839 ? 32'h0/* 0*/ : rb1RowAddr_7;
  assign T1372 = T1380 | T1373;
  assign T1373 = rb1RowAddr_6 & T1374;
  assign T1374 = {6'h20/* 32*/{T764}};
  assign T1375 = T849 || T1376;
  assign T1376 = T1360 && T764;
  assign T1377 = T1376 ? r : T1378;
  assign T1378 = {28'h0/* 0*/, T1379};
  assign T1379 = T849 ? 32'h0/* 0*/ : rb1RowAddr_6;
  assign T1380 = T1387 | T1381;
  assign T1381 = rb1RowAddr_5 & T1382;
  assign T1382 = {6'h20/* 32*/{T777}};
  assign T1383 = T855 || T1359;
  assign T1384 = T1359 ? r : T1385;
  assign T1385 = {28'h0/* 0*/, T1386};
  assign T1386 = T855 ? 32'h0/* 0*/ : rb1RowAddr_5;
  assign T1387 = T1395 | T1388;
  assign T1388 = rb1RowAddr_4 & T1389;
  assign T1389 = {6'h20/* 32*/{T861}};
  assign T1390 = T862 || T1391;
  assign T1391 = T1360 && T861;
  assign T1392 = T1391 ? r : T1393;
  assign T1393 = {28'h0/* 0*/, T1394};
  assign T1394 = T862 ? 32'h0/* 0*/ : rb1RowAddr_4;
  assign T1395 = T1403 | T1396;
  assign T1396 = rb1RowAddr_3 & T1397;
  assign T1397 = {6'h20/* 32*/{T868}};
  assign T1398 = T869 || T1399;
  assign T1399 = T1360 && T868;
  assign T1400 = T1399 ? r : T1401;
  assign T1401 = {28'h0/* 0*/, T1402};
  assign T1402 = T869 ? 32'h0/* 0*/ : rb1RowAddr_3;
  assign T1403 = T1411 | T1404;
  assign T1404 = rb1RowAddr_2 & T1405;
  assign T1405 = {6'h20/* 32*/{T875}};
  assign T1406 = T876 || T1407;
  assign T1407 = T1360 && T875;
  assign T1408 = T1407 ? r : T1409;
  assign T1409 = {28'h0/* 0*/, T1410};
  assign T1410 = T876 ? 32'h0/* 0*/ : rb1RowAddr_2;
  assign T1411 = T1419 | T1412;
  assign T1412 = rb1RowAddr_1 & T1413;
  assign T1413 = {6'h20/* 32*/{T882}};
  assign T1414 = T883 || T1415;
  assign T1415 = T1360 && T882;
  assign T1416 = T1415 ? r : T1417;
  assign T1417 = {28'h0/* 0*/, T1418};
  assign T1418 = T883 ? 32'h0/* 0*/ : rb1RowAddr_1;
  assign T1419 = rb1RowAddr_0 & T1420;
  assign T1420 = {6'h20/* 32*/{T888}};
  assign T1421 = T889 || T1422;
  assign T1422 = T1360 && T888;
  assign T1423 = T1422 ? r : T1424;
  assign T1424 = {28'h0/* 0*/, T1425};
  assign T1425 = T889 ? 32'h0/* 0*/ : rb1RowAddr_0;
  assign T1426 = T916 && T914;
  assign T1427 = T1430 || T1428;
  assign T1428 = T1429 && T777;
  assign T1429 = T1426 && T1362;
  assign T1430 = T1499 || T1431;
  assign T1431 = T1432 && T777;
  assign T1432 = T1498 && T1433;
  assign T1433 = ! T1434;
  assign T1434 = T1435 == r;
  assign T1435 = {28'h0/* 0*/, T1436};
  assign T1436 = T1444 | T1437;
  assign T1437 = rb0RowAddr_7 & T1438;
  assign T1438 = {6'h20/* 32*/{T5}};
  assign T1439 = T839 || T1440;
  assign T1440 = T1432 && T5;
  assign T1441 = T1440 ? r : T1442;
  assign T1442 = {28'h0/* 0*/, T1443};
  assign T1443 = T839 ? 32'h1/* 1*/ : rb0RowAddr_7;
  assign T1444 = T1452 | T1445;
  assign T1445 = rb0RowAddr_6 & T1446;
  assign T1446 = {6'h20/* 32*/{T764}};
  assign T1447 = T849 || T1448;
  assign T1448 = T1432 && T764;
  assign T1449 = T1448 ? r : T1450;
  assign T1450 = {28'h0/* 0*/, T1451};
  assign T1451 = T849 ? 32'h1/* 1*/ : rb0RowAddr_6;
  assign T1452 = T1459 | T1453;
  assign T1453 = rb0RowAddr_5 & T1454;
  assign T1454 = {6'h20/* 32*/{T777}};
  assign T1455 = T855 || T1431;
  assign T1456 = T1431 ? r : T1457;
  assign T1457 = {28'h0/* 0*/, T1458};
  assign T1458 = T855 ? 32'h1/* 1*/ : rb0RowAddr_5;
  assign T1459 = T1467 | T1460;
  assign T1460 = rb0RowAddr_4 & T1461;
  assign T1461 = {6'h20/* 32*/{T861}};
  assign T1462 = T862 || T1463;
  assign T1463 = T1432 && T861;
  assign T1464 = T1463 ? r : T1465;
  assign T1465 = {28'h0/* 0*/, T1466};
  assign T1466 = T862 ? 32'h1/* 1*/ : rb0RowAddr_4;
  assign T1467 = T1475 | T1468;
  assign T1468 = rb0RowAddr_3 & T1469;
  assign T1469 = {6'h20/* 32*/{T868}};
  assign T1470 = T869 || T1471;
  assign T1471 = T1432 && T868;
  assign T1472 = T1471 ? r : T1473;
  assign T1473 = {28'h0/* 0*/, T1474};
  assign T1474 = T869 ? 32'h1/* 1*/ : rb0RowAddr_3;
  assign T1475 = T1483 | T1476;
  assign T1476 = rb0RowAddr_2 & T1477;
  assign T1477 = {6'h20/* 32*/{T875}};
  assign T1478 = T876 || T1479;
  assign T1479 = T1432 && T875;
  assign T1480 = T1479 ? r : T1481;
  assign T1481 = {28'h0/* 0*/, T1482};
  assign T1482 = T876 ? 32'h1/* 1*/ : rb0RowAddr_2;
  assign T1483 = T1491 | T1484;
  assign T1484 = rb0RowAddr_1 & T1485;
  assign T1485 = {6'h20/* 32*/{T882}};
  assign T1486 = T883 || T1487;
  assign T1487 = T1432 && T882;
  assign T1488 = T1487 ? r : T1489;
  assign T1489 = {28'h0/* 0*/, T1490};
  assign T1490 = T883 ? 32'h1/* 1*/ : rb0RowAddr_1;
  assign T1491 = rb0RowAddr_0 & T1492;
  assign T1492 = {6'h20/* 32*/{T888}};
  assign T1493 = T889 || T1494;
  assign T1494 = T1432 && T888;
  assign T1495 = T1494 ? r : T1496;
  assign T1496 = {28'h0/* 0*/, T1497};
  assign T1497 = T889 ? 32'h1/* 1*/ : rb0RowAddr_0;
  assign T1498 = T920 && T918;
  assign T1499 = T1502 || T1500;
  assign T1500 = T1501 && T777;
  assign T1501 = T1498 && T1434;
  assign T1502 = T855 || T1503;
  assign T1503 = T1504 && T84;
  assign T1504 = T1505 && io_out_ready;
  assign T1505 = T1507 && T1506;
  assign T1506 = T19 == 8'hff/* 255*/;
  assign T1507 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T1508 = T1766 ? 8'hff/* 255*/ : T1509;
  assign T1509 = T829 ? T1765 : T1510;
  assign T1510 = T925 ? T1764 : T1511;
  assign T1511 = T996 ? T1763 : T1512;
  assign T1512 = T999 ? T1762 : T1513;
  assign T1513 = T1068 ? T1761 : T1514;
  assign T1514 = T1071 ? T1760 : T1515;
  assign T1515 = T1140 ? T1759 : T1516;
  assign T1516 = T1143 ? T1758 : T1517;
  assign T1517 = T1212 ? T1757 : T1518;
  assign T1518 = T1215 ? T1756 : T1519;
  assign T1519 = T1284 ? T1755 : T1520;
  assign T1520 = T1287 ? T1754 : T1521;
  assign T1521 = T1356 ? T1753 : T1522;
  assign T1522 = T1359 ? T1752 : T1523;
  assign T1523 = T1428 ? T1751 : T1524;
  assign T1524 = T1431 ? T1750 : T1525;
  assign T1525 = T1500 ? T1749 : T1526;
  assign T1526 = T1503 ? T1529 : T1527;
  assign T1527 = T855 ? T1528 : State_5;
  assign T1528 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1529 = T1557 | T1530;
  assign T1530 = EmitReturnState_7 & T1531;
  assign T1531 = {4'h8/* 8*/{T22}};
  assign T1532 = T1533 || T4;
  assign T1533 = T1535 || T1534;
  assign T1534 = T782 && T5;
  assign T1535 = T1537 || T1536;
  assign T1536 = T788 && T5;
  assign T1537 = T1539 || T1538;
  assign T1538 = T794 && T5;
  assign T1539 = T1541 || T1540;
  assign T1540 = T800 && T5;
  assign T1541 = T1543 || T1542;
  assign T1542 = T806 && T5;
  assign T1543 = T1545 || T1544;
  assign T1544 = T812 && T5;
  assign T1545 = T1547 || T1546;
  assign T1546 = T818 && T5;
  assign T1547 = T824 && T5;
  assign T1548 = T1549 ? 8'h0/* 0*/ : EmitReturnState_7;
  assign T1549 = T1550 || T4;
  assign T1550 = T1551 || T1534;
  assign T1551 = T1552 || T1536;
  assign T1552 = T1553 || T1538;
  assign T1553 = T1554 || T1540;
  assign T1554 = T1555 || T1542;
  assign T1555 = T1556 || T1544;
  assign T1556 = T1547 || T1546;
  assign T1557 = T1585 | T1558;
  assign T1558 = EmitReturnState_6 & T1559;
  assign T1559 = {4'h8/* 8*/{T73}};
  assign T1560 = T1561 || T763;
  assign T1561 = T1563 || T1562;
  assign T1562 = T782 && T764;
  assign T1563 = T1565 || T1564;
  assign T1564 = T788 && T764;
  assign T1565 = T1567 || T1566;
  assign T1566 = T794 && T764;
  assign T1567 = T1569 || T1568;
  assign T1568 = T800 && T764;
  assign T1569 = T1571 || T1570;
  assign T1570 = T806 && T764;
  assign T1571 = T1573 || T1572;
  assign T1572 = T812 && T764;
  assign T1573 = T1575 || T1574;
  assign T1574 = T818 && T764;
  assign T1575 = T824 && T764;
  assign T1576 = T1577 ? 8'h0/* 0*/ : EmitReturnState_6;
  assign T1577 = T1578 || T763;
  assign T1578 = T1579 || T1562;
  assign T1579 = T1580 || T1564;
  assign T1580 = T1581 || T1566;
  assign T1581 = T1582 || T1568;
  assign T1582 = T1583 || T1570;
  assign T1583 = T1584 || T1572;
  assign T1584 = T1575 || T1574;
  assign T1585 = T1605 | T1586;
  assign T1586 = EmitReturnState_5 & T1587;
  assign T1587 = {4'h8/* 8*/{T84}};
  assign T1588 = T1589 || T779;
  assign T1589 = T1590 || T781;
  assign T1590 = T1591 || T787;
  assign T1591 = T1592 || T793;
  assign T1592 = T1593 || T799;
  assign T1593 = T1594 || T805;
  assign T1594 = T1595 || T811;
  assign T1595 = T823 || T817;
  assign T1596 = T1597 ? 8'h0/* 0*/ : EmitReturnState_5;
  assign T1597 = T1598 || T779;
  assign T1598 = T1599 || T781;
  assign T1599 = T1600 || T787;
  assign T1600 = T1601 || T793;
  assign T1601 = T1602 || T799;
  assign T1602 = T1603 || T805;
  assign T1603 = T1604 || T811;
  assign T1604 = T823 || T817;
  assign T1605 = T1634 | T1606;
  assign T1606 = EmitReturnState_4 & T1607;
  assign T1607 = {4'h8/* 8*/{T95}};
  assign T1608 = T1610 || T1609;
  assign T1609 = T765 && T861;
  assign T1610 = T1612 || T1611;
  assign T1611 = T782 && T861;
  assign T1612 = T1614 || T1613;
  assign T1613 = T788 && T861;
  assign T1614 = T1616 || T1615;
  assign T1615 = T794 && T861;
  assign T1616 = T1618 || T1617;
  assign T1617 = T800 && T861;
  assign T1618 = T1620 || T1619;
  assign T1619 = T806 && T861;
  assign T1620 = T1622 || T1621;
  assign T1621 = T812 && T861;
  assign T1622 = T1624 || T1623;
  assign T1623 = T818 && T861;
  assign T1624 = T824 && T861;
  assign T1625 = T1626 ? 8'h0/* 0*/ : EmitReturnState_4;
  assign T1626 = T1627 || T1609;
  assign T1627 = T1628 || T1611;
  assign T1628 = T1629 || T1613;
  assign T1629 = T1630 || T1615;
  assign T1630 = T1631 || T1617;
  assign T1631 = T1632 || T1619;
  assign T1632 = T1633 || T1621;
  assign T1633 = T1624 || T1623;
  assign T1634 = T1663 | T1635;
  assign T1635 = EmitReturnState_3 & T1636;
  assign T1636 = {4'h8/* 8*/{T106}};
  assign T1637 = T1639 || T1638;
  assign T1638 = T765 && T868;
  assign T1639 = T1641 || T1640;
  assign T1640 = T782 && T868;
  assign T1641 = T1643 || T1642;
  assign T1642 = T788 && T868;
  assign T1643 = T1645 || T1644;
  assign T1644 = T794 && T868;
  assign T1645 = T1647 || T1646;
  assign T1646 = T800 && T868;
  assign T1647 = T1649 || T1648;
  assign T1648 = T806 && T868;
  assign T1649 = T1651 || T1650;
  assign T1650 = T812 && T868;
  assign T1651 = T1653 || T1652;
  assign T1652 = T818 && T868;
  assign T1653 = T824 && T868;
  assign T1654 = T1655 ? 8'h0/* 0*/ : EmitReturnState_3;
  assign T1655 = T1656 || T1638;
  assign T1656 = T1657 || T1640;
  assign T1657 = T1658 || T1642;
  assign T1658 = T1659 || T1644;
  assign T1659 = T1660 || T1646;
  assign T1660 = T1661 || T1648;
  assign T1661 = T1662 || T1650;
  assign T1662 = T1653 || T1652;
  assign T1663 = T1692 | T1664;
  assign T1664 = EmitReturnState_2 & T1665;
  assign T1665 = {4'h8/* 8*/{T117}};
  assign T1666 = T1668 || T1667;
  assign T1667 = T765 && T875;
  assign T1668 = T1670 || T1669;
  assign T1669 = T782 && T875;
  assign T1670 = T1672 || T1671;
  assign T1671 = T788 && T875;
  assign T1672 = T1674 || T1673;
  assign T1673 = T794 && T875;
  assign T1674 = T1676 || T1675;
  assign T1675 = T800 && T875;
  assign T1676 = T1678 || T1677;
  assign T1677 = T806 && T875;
  assign T1678 = T1680 || T1679;
  assign T1679 = T812 && T875;
  assign T1680 = T1682 || T1681;
  assign T1681 = T818 && T875;
  assign T1682 = T824 && T875;
  assign T1683 = T1684 ? 8'h0/* 0*/ : EmitReturnState_2;
  assign T1684 = T1685 || T1667;
  assign T1685 = T1686 || T1669;
  assign T1686 = T1687 || T1671;
  assign T1687 = T1688 || T1673;
  assign T1688 = T1689 || T1675;
  assign T1689 = T1690 || T1677;
  assign T1690 = T1691 || T1679;
  assign T1691 = T1682 || T1681;
  assign T1692 = T1721 | T1693;
  assign T1693 = EmitReturnState_1 & T1694;
  assign T1694 = {4'h8/* 8*/{T128}};
  assign T1695 = T1697 || T1696;
  assign T1696 = T765 && T882;
  assign T1697 = T1699 || T1698;
  assign T1698 = T782 && T882;
  assign T1699 = T1701 || T1700;
  assign T1700 = T788 && T882;
  assign T1701 = T1703 || T1702;
  assign T1702 = T794 && T882;
  assign T1703 = T1705 || T1704;
  assign T1704 = T800 && T882;
  assign T1705 = T1707 || T1706;
  assign T1706 = T806 && T882;
  assign T1707 = T1709 || T1708;
  assign T1708 = T812 && T882;
  assign T1709 = T1711 || T1710;
  assign T1710 = T818 && T882;
  assign T1711 = T824 && T882;
  assign T1712 = T1713 ? 8'h0/* 0*/ : EmitReturnState_1;
  assign T1713 = T1714 || T1696;
  assign T1714 = T1715 || T1698;
  assign T1715 = T1716 || T1700;
  assign T1716 = T1717 || T1702;
  assign T1717 = T1718 || T1704;
  assign T1718 = T1719 || T1706;
  assign T1719 = T1720 || T1708;
  assign T1720 = T1711 || T1710;
  assign T1721 = EmitReturnState_0 & T1722;
  assign T1722 = {4'h8/* 8*/{T138}};
  assign T1723 = T1725 || T1724;
  assign T1724 = T765 && T888;
  assign T1725 = T1727 || T1726;
  assign T1726 = T782 && T888;
  assign T1727 = T1729 || T1728;
  assign T1728 = T788 && T888;
  assign T1729 = T1731 || T1730;
  assign T1730 = T794 && T888;
  assign T1731 = T1733 || T1732;
  assign T1732 = T800 && T888;
  assign T1733 = T1735 || T1734;
  assign T1734 = T806 && T888;
  assign T1735 = T1737 || T1736;
  assign T1736 = T812 && T888;
  assign T1737 = T1739 || T1738;
  assign T1738 = T818 && T888;
  assign T1739 = T824 && T888;
  assign T1740 = T1741 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T1741 = T1742 || T1724;
  assign T1742 = T1743 || T1726;
  assign T1743 = T1744 || T1728;
  assign T1744 = T1745 || T1730;
  assign T1745 = T1746 || T1732;
  assign T1746 = T1747 || T1734;
  assign T1747 = T1748 || T1736;
  assign T1748 = T1739 || T1738;
  assign T1749 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1750 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1751 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1752 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1753 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1754 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1755 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1756 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1757 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1758 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1759 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1760 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1761 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1762 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1763 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1764 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1765 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1766 = T1767 || T779;
  assign T1767 = T1768 || T781;
  assign T1768 = T1769 || T787;
  assign T1769 = T1770 || T793;
  assign T1770 = T1771 || T799;
  assign T1771 = T1772 || T805;
  assign T1772 = T1773 || T811;
  assign T1773 = T823 || T817;
  assign T1774 = T1860 | T1775;
  assign T1775 = State_4 & T1776;
  assign T1776 = {4'h8/* 8*/{T861}};
  assign T1777 = T1778 || T1609;
  assign T1778 = T1779 || T1611;
  assign T1779 = T1780 || T1613;
  assign T1780 = T1781 || T1615;
  assign T1781 = T1782 || T1617;
  assign T1782 = T1783 || T1619;
  assign T1783 = T1784 || T1621;
  assign T1784 = T1785 || T1623;
  assign T1785 = T1786 || T1624;
  assign T1786 = T1788 || T1787;
  assign T1787 = T830 && T861;
  assign T1788 = T1789 || T959;
  assign T1789 = T1791 || T1790;
  assign T1790 = T997 && T861;
  assign T1791 = T1792 || T1031;
  assign T1792 = T1794 || T1793;
  assign T1793 = T1069 && T861;
  assign T1794 = T1795 || T1103;
  assign T1795 = T1797 || T1796;
  assign T1796 = T1141 && T861;
  assign T1797 = T1798 || T1175;
  assign T1798 = T1800 || T1799;
  assign T1799 = T1213 && T861;
  assign T1800 = T1801 || T1247;
  assign T1801 = T1803 || T1802;
  assign T1802 = T1285 && T861;
  assign T1803 = T1804 || T1319;
  assign T1804 = T1806 || T1805;
  assign T1805 = T1357 && T861;
  assign T1806 = T1807 || T1391;
  assign T1807 = T1809 || T1808;
  assign T1808 = T1429 && T861;
  assign T1809 = T1810 || T1463;
  assign T1810 = T1812 || T1811;
  assign T1811 = T1501 && T861;
  assign T1812 = T862 || T1813;
  assign T1813 = T1504 && T95;
  assign T1814 = T1852 ? 8'hff/* 255*/ : T1815;
  assign T1815 = T1787 ? T1851 : T1816;
  assign T1816 = T959 ? T1850 : T1817;
  assign T1817 = T1790 ? T1849 : T1818;
  assign T1818 = T1031 ? T1848 : T1819;
  assign T1819 = T1793 ? T1847 : T1820;
  assign T1820 = T1103 ? T1846 : T1821;
  assign T1821 = T1796 ? T1845 : T1822;
  assign T1822 = T1175 ? T1844 : T1823;
  assign T1823 = T1799 ? T1843 : T1824;
  assign T1824 = T1247 ? T1842 : T1825;
  assign T1825 = T1802 ? T1841 : T1826;
  assign T1826 = T1319 ? T1840 : T1827;
  assign T1827 = T1805 ? T1839 : T1828;
  assign T1828 = T1391 ? T1838 : T1829;
  assign T1829 = T1808 ? T1837 : T1830;
  assign T1830 = T1463 ? T1836 : T1831;
  assign T1831 = T1811 ? T1835 : T1832;
  assign T1832 = T1813 ? T1529 : T1833;
  assign T1833 = T862 ? T1834 : State_4;
  assign T1834 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1835 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1836 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1837 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1838 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1839 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1840 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1841 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1842 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1843 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1844 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1845 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1846 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1847 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1848 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1849 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1850 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1851 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1852 = T1853 || T1609;
  assign T1853 = T1854 || T1611;
  assign T1854 = T1855 || T1613;
  assign T1855 = T1856 || T1615;
  assign T1856 = T1857 || T1617;
  assign T1857 = T1858 || T1619;
  assign T1858 = T1859 || T1621;
  assign T1859 = T1624 || T1623;
  assign T1860 = T1946 | T1861;
  assign T1861 = State_3 & T1862;
  assign T1862 = {4'h8/* 8*/{T868}};
  assign T1863 = T1864 || T1638;
  assign T1864 = T1865 || T1640;
  assign T1865 = T1866 || T1642;
  assign T1866 = T1867 || T1644;
  assign T1867 = T1868 || T1646;
  assign T1868 = T1869 || T1648;
  assign T1869 = T1870 || T1650;
  assign T1870 = T1871 || T1652;
  assign T1871 = T1872 || T1653;
  assign T1872 = T1874 || T1873;
  assign T1873 = T830 && T868;
  assign T1874 = T1875 || T967;
  assign T1875 = T1877 || T1876;
  assign T1876 = T997 && T868;
  assign T1877 = T1878 || T1039;
  assign T1878 = T1880 || T1879;
  assign T1879 = T1069 && T868;
  assign T1880 = T1881 || T1111;
  assign T1881 = T1883 || T1882;
  assign T1882 = T1141 && T868;
  assign T1883 = T1884 || T1183;
  assign T1884 = T1886 || T1885;
  assign T1885 = T1213 && T868;
  assign T1886 = T1887 || T1255;
  assign T1887 = T1889 || T1888;
  assign T1888 = T1285 && T868;
  assign T1889 = T1890 || T1327;
  assign T1890 = T1892 || T1891;
  assign T1891 = T1357 && T868;
  assign T1892 = T1893 || T1399;
  assign T1893 = T1895 || T1894;
  assign T1894 = T1429 && T868;
  assign T1895 = T1896 || T1471;
  assign T1896 = T1898 || T1897;
  assign T1897 = T1501 && T868;
  assign T1898 = T869 || T1899;
  assign T1899 = T1504 && T106;
  assign T1900 = T1938 ? 8'hff/* 255*/ : T1901;
  assign T1901 = T1873 ? T1937 : T1902;
  assign T1902 = T967 ? T1936 : T1903;
  assign T1903 = T1876 ? T1935 : T1904;
  assign T1904 = T1039 ? T1934 : T1905;
  assign T1905 = T1879 ? T1933 : T1906;
  assign T1906 = T1111 ? T1932 : T1907;
  assign T1907 = T1882 ? T1931 : T1908;
  assign T1908 = T1183 ? T1930 : T1909;
  assign T1909 = T1885 ? T1929 : T1910;
  assign T1910 = T1255 ? T1928 : T1911;
  assign T1911 = T1888 ? T1927 : T1912;
  assign T1912 = T1327 ? T1926 : T1913;
  assign T1913 = T1891 ? T1925 : T1914;
  assign T1914 = T1399 ? T1924 : T1915;
  assign T1915 = T1894 ? T1923 : T1916;
  assign T1916 = T1471 ? T1922 : T1917;
  assign T1917 = T1897 ? T1921 : T1918;
  assign T1918 = T1899 ? T1529 : T1919;
  assign T1919 = T869 ? T1920 : State_3;
  assign T1920 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T1921 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1922 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T1923 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1924 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T1925 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1926 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T1927 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1928 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T1929 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1930 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T1931 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1932 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T1933 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1934 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T1935 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1936 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T1937 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T1938 = T1939 || T1638;
  assign T1939 = T1940 || T1640;
  assign T1940 = T1941 || T1642;
  assign T1941 = T1942 || T1644;
  assign T1942 = T1943 || T1646;
  assign T1943 = T1944 || T1648;
  assign T1944 = T1945 || T1650;
  assign T1945 = T1653 || T1652;
  assign T1946 = T2032 | T1947;
  assign T1947 = State_2 & T1948;
  assign T1948 = {4'h8/* 8*/{T875}};
  assign T1949 = T1950 || T1667;
  assign T1950 = T1951 || T1669;
  assign T1951 = T1952 || T1671;
  assign T1952 = T1953 || T1673;
  assign T1953 = T1954 || T1675;
  assign T1954 = T1955 || T1677;
  assign T1955 = T1956 || T1679;
  assign T1956 = T1957 || T1681;
  assign T1957 = T1958 || T1682;
  assign T1958 = T1960 || T1959;
  assign T1959 = T830 && T875;
  assign T1960 = T1961 || T975;
  assign T1961 = T1963 || T1962;
  assign T1962 = T997 && T875;
  assign T1963 = T1964 || T1047;
  assign T1964 = T1966 || T1965;
  assign T1965 = T1069 && T875;
  assign T1966 = T1967 || T1119;
  assign T1967 = T1969 || T1968;
  assign T1968 = T1141 && T875;
  assign T1969 = T1970 || T1191;
  assign T1970 = T1972 || T1971;
  assign T1971 = T1213 && T875;
  assign T1972 = T1973 || T1263;
  assign T1973 = T1975 || T1974;
  assign T1974 = T1285 && T875;
  assign T1975 = T1976 || T1335;
  assign T1976 = T1978 || T1977;
  assign T1977 = T1357 && T875;
  assign T1978 = T1979 || T1407;
  assign T1979 = T1981 || T1980;
  assign T1980 = T1429 && T875;
  assign T1981 = T1982 || T1479;
  assign T1982 = T1984 || T1983;
  assign T1983 = T1501 && T875;
  assign T1984 = T876 || T1985;
  assign T1985 = T1504 && T117;
  assign T1986 = T2024 ? 8'hff/* 255*/ : T1987;
  assign T1987 = T1959 ? T2023 : T1988;
  assign T1988 = T975 ? T2022 : T1989;
  assign T1989 = T1962 ? T2021 : T1990;
  assign T1990 = T1047 ? T2020 : T1991;
  assign T1991 = T1965 ? T2019 : T1992;
  assign T1992 = T1119 ? T2018 : T1993;
  assign T1993 = T1968 ? T2017 : T1994;
  assign T1994 = T1191 ? T2016 : T1995;
  assign T1995 = T1971 ? T2015 : T1996;
  assign T1996 = T1263 ? T2014 : T1997;
  assign T1997 = T1974 ? T2013 : T1998;
  assign T1998 = T1335 ? T2012 : T1999;
  assign T1999 = T1977 ? T2011 : T2000;
  assign T2000 = T1407 ? T2010 : T2001;
  assign T2001 = T1980 ? T2009 : T2002;
  assign T2002 = T1479 ? T2008 : T2003;
  assign T2003 = T1983 ? T2007 : T2004;
  assign T2004 = T1985 ? T1529 : T2005;
  assign T2005 = T876 ? T2006 : State_2;
  assign T2006 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2007 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2008 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2009 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2010 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2011 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2012 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2013 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2014 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2015 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2016 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2017 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2018 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2019 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2020 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2021 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2022 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2023 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2024 = T2025 || T1667;
  assign T2025 = T2026 || T1669;
  assign T2026 = T2027 || T1671;
  assign T2027 = T2028 || T1673;
  assign T2028 = T2029 || T1675;
  assign T2029 = T2030 || T1677;
  assign T2030 = T2031 || T1679;
  assign T2031 = T1682 || T1681;
  assign T2032 = T2118 | T2033;
  assign T2033 = State_1 & T2034;
  assign T2034 = {4'h8/* 8*/{T882}};
  assign T2035 = T2036 || T1696;
  assign T2036 = T2037 || T1698;
  assign T2037 = T2038 || T1700;
  assign T2038 = T2039 || T1702;
  assign T2039 = T2040 || T1704;
  assign T2040 = T2041 || T1706;
  assign T2041 = T2042 || T1708;
  assign T2042 = T2043 || T1710;
  assign T2043 = T2044 || T1711;
  assign T2044 = T2046 || T2045;
  assign T2045 = T830 && T882;
  assign T2046 = T2047 || T983;
  assign T2047 = T2049 || T2048;
  assign T2048 = T997 && T882;
  assign T2049 = T2050 || T1055;
  assign T2050 = T2052 || T2051;
  assign T2051 = T1069 && T882;
  assign T2052 = T2053 || T1127;
  assign T2053 = T2055 || T2054;
  assign T2054 = T1141 && T882;
  assign T2055 = T2056 || T1199;
  assign T2056 = T2058 || T2057;
  assign T2057 = T1213 && T882;
  assign T2058 = T2059 || T1271;
  assign T2059 = T2061 || T2060;
  assign T2060 = T1285 && T882;
  assign T2061 = T2062 || T1343;
  assign T2062 = T2064 || T2063;
  assign T2063 = T1357 && T882;
  assign T2064 = T2065 || T1415;
  assign T2065 = T2067 || T2066;
  assign T2066 = T1429 && T882;
  assign T2067 = T2068 || T1487;
  assign T2068 = T2070 || T2069;
  assign T2069 = T1501 && T882;
  assign T2070 = T883 || T2071;
  assign T2071 = T1504 && T128;
  assign T2072 = T2110 ? 8'hff/* 255*/ : T2073;
  assign T2073 = T2045 ? T2109 : T2074;
  assign T2074 = T983 ? T2108 : T2075;
  assign T2075 = T2048 ? T2107 : T2076;
  assign T2076 = T1055 ? T2106 : T2077;
  assign T2077 = T2051 ? T2105 : T2078;
  assign T2078 = T1127 ? T2104 : T2079;
  assign T2079 = T2054 ? T2103 : T2080;
  assign T2080 = T1199 ? T2102 : T2081;
  assign T2081 = T2057 ? T2101 : T2082;
  assign T2082 = T1271 ? T2100 : T2083;
  assign T2083 = T2060 ? T2099 : T2084;
  assign T2084 = T1343 ? T2098 : T2085;
  assign T2085 = T2063 ? T2097 : T2086;
  assign T2086 = T1415 ? T2096 : T2087;
  assign T2087 = T2066 ? T2095 : T2088;
  assign T2088 = T1487 ? T2094 : T2089;
  assign T2089 = T2069 ? T2093 : T2090;
  assign T2090 = T2071 ? T1529 : T2091;
  assign T2091 = T883 ? T2092 : State_1;
  assign T2092 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2093 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2094 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2095 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2096 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2097 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2098 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2099 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2100 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2101 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2102 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2103 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2104 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2105 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2106 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2107 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2108 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2109 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2110 = T2111 || T1696;
  assign T2111 = T2112 || T1698;
  assign T2112 = T2113 || T1700;
  assign T2113 = T2114 || T1702;
  assign T2114 = T2115 || T1704;
  assign T2115 = T2116 || T1706;
  assign T2116 = T2117 || T1708;
  assign T2117 = T1711 || T1710;
  assign T2118 = State_0 & T2119;
  assign T2119 = {4'h8/* 8*/{T888}};
  assign T2120 = T2121 || T1724;
  assign T2121 = T2122 || T1726;
  assign T2122 = T2123 || T1728;
  assign T2123 = T2124 || T1730;
  assign T2124 = T2125 || T1732;
  assign T2125 = T2126 || T1734;
  assign T2126 = T2127 || T1736;
  assign T2127 = T2128 || T1738;
  assign T2128 = T2129 || T1739;
  assign T2129 = T2131 || T2130;
  assign T2130 = T830 && T888;
  assign T2131 = T2132 || T990;
  assign T2132 = T2134 || T2133;
  assign T2133 = T997 && T888;
  assign T2134 = T2135 || T1062;
  assign T2135 = T2137 || T2136;
  assign T2136 = T1069 && T888;
  assign T2137 = T2138 || T1134;
  assign T2138 = T2140 || T2139;
  assign T2139 = T1141 && T888;
  assign T2140 = T2141 || T1206;
  assign T2141 = T2143 || T2142;
  assign T2142 = T1213 && T888;
  assign T2143 = T2144 || T1278;
  assign T2144 = T2146 || T2145;
  assign T2145 = T1285 && T888;
  assign T2146 = T2147 || T1350;
  assign T2147 = T2149 || T2148;
  assign T2148 = T1357 && T888;
  assign T2149 = T2150 || T1422;
  assign T2150 = T2152 || T2151;
  assign T2151 = T1429 && T888;
  assign T2152 = T2153 || T1494;
  assign T2153 = T2155 || T2154;
  assign T2154 = T1501 && T888;
  assign T2155 = T889 || T2156;
  assign T2156 = T1504 && T138;
  assign T2157 = T2195 ? 8'hff/* 255*/ : T2158;
  assign T2158 = T2130 ? T2194 : T2159;
  assign T2159 = T990 ? T2193 : T2160;
  assign T2160 = T2133 ? T2192 : T2161;
  assign T2161 = T1062 ? T2191 : T2162;
  assign T2162 = T2136 ? T2190 : T2163;
  assign T2163 = T1134 ? T2189 : T2164;
  assign T2164 = T2139 ? T2188 : T2165;
  assign T2165 = T1206 ? T2187 : T2166;
  assign T2166 = T2142 ? T2186 : T2167;
  assign T2167 = T1278 ? T2185 : T2168;
  assign T2168 = T2145 ? T2184 : T2169;
  assign T2169 = T1350 ? T2183 : T2170;
  assign T2170 = T2148 ? T2182 : T2171;
  assign T2171 = T1422 ? T2181 : T2172;
  assign T2172 = T2151 ? T2180 : T2173;
  assign T2173 = T1494 ? T2179 : T2174;
  assign T2174 = T2154 ? T2178 : T2175;
  assign T2175 = T2156 ? T1529 : T2176;
  assign T2176 = T889 ? T2177 : State_0;
  assign T2177 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2178 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2179 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2180 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2181 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2182 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2183 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2184 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2185 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2186 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2187 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2188 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2189 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2190 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2191 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2192 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2193 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2194 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2195 = T2196 || T1724;
  assign T2196 = T2197 || T1726;
  assign T2197 = T2198 || T1728;
  assign T2198 = T2199 || T1730;
  assign T2199 = T2200 || T1732;
  assign T2200 = T2201 || T1734;
  assign T2201 = T2202 || T1736;
  assign T2202 = T1739 || T1738;
  assign T2203 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2204 = T2205 || T1562;
  assign T2205 = T2206 || T1564;
  assign T2206 = T2207 || T1566;
  assign T2207 = T2208 || T1568;
  assign T2208 = T2209 || T1570;
  assign T2209 = T2210 || T1572;
  assign T2210 = T2211 || T1574;
  assign T2211 = T2212 || T1575;
  assign T2212 = T2214 || T2213;
  assign T2213 = T830 && T764;
  assign T2214 = T2215 || T944;
  assign T2215 = T2217 || T2216;
  assign T2216 = T997 && T764;
  assign T2217 = T2218 || T1016;
  assign T2218 = T2220 || T2219;
  assign T2219 = T1069 && T764;
  assign T2220 = T2221 || T1088;
  assign T2221 = T2223 || T2222;
  assign T2222 = T1141 && T764;
  assign T2223 = T2224 || T1160;
  assign T2224 = T2226 || T2225;
  assign T2225 = T1213 && T764;
  assign T2226 = T2227 || T1232;
  assign T2227 = T2229 || T2228;
  assign T2228 = T1285 && T764;
  assign T2229 = T2230 || T1304;
  assign T2230 = T2232 || T2231;
  assign T2231 = T1357 && T764;
  assign T2232 = T2233 || T1376;
  assign T2233 = T2235 || T2234;
  assign T2234 = T1429 && T764;
  assign T2235 = T2236 || T1448;
  assign T2236 = T2238 || T2237;
  assign T2237 = T1501 && T764;
  assign T2238 = T849 || T2239;
  assign T2239 = T1504 && T73;
  assign T2240 = T2278 ? 8'hff/* 255*/ : T2241;
  assign T2241 = T2213 ? T2277 : T2242;
  assign T2242 = T944 ? T2276 : T2243;
  assign T2243 = T2216 ? T2275 : T2244;
  assign T2244 = T1016 ? T2274 : T2245;
  assign T2245 = T2219 ? T2273 : T2246;
  assign T2246 = T1088 ? T2272 : T2247;
  assign T2247 = T2222 ? T2271 : T2248;
  assign T2248 = T1160 ? T2270 : T2249;
  assign T2249 = T2225 ? T2269 : T2250;
  assign T2250 = T1232 ? T2268 : T2251;
  assign T2251 = T2228 ? T2267 : T2252;
  assign T2252 = T1304 ? T2266 : T2253;
  assign T2253 = T2231 ? T2265 : T2254;
  assign T2254 = T1376 ? T2264 : T2255;
  assign T2255 = T2234 ? T2263 : T2256;
  assign T2256 = T1448 ? T2262 : T2257;
  assign T2257 = T2237 ? T2261 : T2258;
  assign T2258 = T2239 ? T1529 : T2259;
  assign T2259 = T849 ? T2260 : State_6;
  assign T2260 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T2261 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2262 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T2263 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2264 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T2265 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2266 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T2267 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2268 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T2269 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2270 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T2271 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2272 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T2273 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2274 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T2275 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2276 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T2277 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T2278 = T2279 || T763;
  assign T2279 = T2280 || T1562;
  assign T2280 = T2281 || T1564;
  assign T2281 = T2282 || T1566;
  assign T2282 = T2283 || T1568;
  assign T2283 = T2284 || T1570;
  assign T2284 = T2285 || T1572;
  assign T2285 = T1575 || T1574;
  assign T2286 = T2288 && T2287;
  assign T2287 = State_6 != 8'h0/* 0*/;
  assign T2288 = AllOffloadsReady && T2289;
  assign T2289 = T2290 == rThreadEncoder_io_chosen;
  assign T2290 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T2291 = subStateTh_5 == 1'h0/* 0*/;
  assign T2292 = T2296 ? 1'h1/* 1*/ : T2293;
  assign T2293 = T2294 ? 1'h0/* 0*/ : subStateTh_5;
  assign T2294 = T2295 == vThreadEncoder_io_chosen;
  assign T2295 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T2296 = T2298 && T2297;
  assign T2297 = State_5 != 8'hff/* 255*/;
  assign T2298 = T2300 && T2299;
  assign T2299 = State_5 != 8'h0/* 0*/;
  assign T2300 = AllOffloadsReady && T2301;
  assign T2301 = T2302 == rThreadEncoder_io_chosen;
  assign T2302 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T2303 = subStateTh_4 == 1'h0/* 0*/;
  assign T2304 = T2308 ? 1'h1/* 1*/ : T2305;
  assign T2305 = T2306 ? 1'h0/* 0*/ : subStateTh_4;
  assign T2306 = T2307 == vThreadEncoder_io_chosen;
  assign T2307 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T2308 = T2310 && T2309;
  assign T2309 = State_4 != 8'hff/* 255*/;
  assign T2310 = T2312 && T2311;
  assign T2311 = State_4 != 8'h0/* 0*/;
  assign T2312 = AllOffloadsReady && T2313;
  assign T2313 = T2314 == rThreadEncoder_io_chosen;
  assign T2314 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T2315 = subStateTh_3 == 1'h0/* 0*/;
  assign T2316 = T2320 ? 1'h1/* 1*/ : T2317;
  assign T2317 = T2318 ? 1'h0/* 0*/ : subStateTh_3;
  assign T2318 = T2319 == vThreadEncoder_io_chosen;
  assign T2319 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T2320 = T2322 && T2321;
  assign T2321 = State_3 != 8'hff/* 255*/;
  assign T2322 = T2324 && T2323;
  assign T2323 = State_3 != 8'h0/* 0*/;
  assign T2324 = AllOffloadsReady && T2325;
  assign T2325 = T2326 == rThreadEncoder_io_chosen;
  assign T2326 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T2327 = subStateTh_2 == 1'h0/* 0*/;
  assign T2328 = T2332 ? 1'h1/* 1*/ : T2329;
  assign T2329 = T2330 ? 1'h0/* 0*/ : subStateTh_2;
  assign T2330 = T2331 == vThreadEncoder_io_chosen;
  assign T2331 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T2332 = T2334 && T2333;
  assign T2333 = State_2 != 8'hff/* 255*/;
  assign T2334 = T2336 && T2335;
  assign T2335 = State_2 != 8'h0/* 0*/;
  assign T2336 = AllOffloadsReady && T2337;
  assign T2337 = T2338 == rThreadEncoder_io_chosen;
  assign T2338 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T2339 = subStateTh_1 == 1'h0/* 0*/;
  assign T2340 = T2344 ? 1'h1/* 1*/ : T2341;
  assign T2341 = T2342 ? 1'h0/* 0*/ : subStateTh_1;
  assign T2342 = T2343 == vThreadEncoder_io_chosen;
  assign T2343 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T2344 = T2346 && T2345;
  assign T2345 = State_1 != 8'hff/* 255*/;
  assign T2346 = T2348 && T2347;
  assign T2347 = State_1 != 8'h0/* 0*/;
  assign T2348 = AllOffloadsReady && T2349;
  assign T2349 = T2350 == rThreadEncoder_io_chosen;
  assign T2350 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T2351 = subStateTh_0 == 1'h0/* 0*/;
  assign T2352 = T2356 ? 1'h1/* 1*/ : T2353;
  assign T2353 = T2354 ? 1'h0/* 0*/ : subStateTh_0;
  assign T2354 = T2355 == vThreadEncoder_io_chosen;
  assign T2355 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T2356 = T2358 && T2357;
  assign T2357 = State_0 != 8'hff/* 255*/;
  assign T2358 = T2360 && T2359;
  assign T2359 = State_0 != 8'h0/* 0*/;
  assign T2360 = AllOffloadsReady && T2361;
  assign T2361 = T2362 == rThreadEncoder_io_chosen;
  assign T2362 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T2363 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2364 = T2367 | T2365;
  assign T2365 = State_6 & T2366;
  assign T2366 = {4'h8/* 8*/{T73}};
  assign T2367 = T2370 | T2368;
  assign T2368 = State_5 & T2369;
  assign T2369 = {4'h8/* 8*/{T84}};
  assign T2370 = T2373 | T2371;
  assign T2371 = State_4 & T2372;
  assign T2372 = {4'h8/* 8*/{T95}};
  assign T2373 = T2376 | T2374;
  assign T2374 = State_3 & T2375;
  assign T2375 = {4'h8/* 8*/{T106}};
  assign T2376 = T2379 | T2377;
  assign T2377 = State_2 & T2378;
  assign T2378 = {4'h8/* 8*/{T117}};
  assign T2379 = T2382 | T2380;
  assign T2380 = State_1 & T2381;
  assign T2381 = {4'h8/* 8*/{T128}};
  assign T2382 = State_0 & T2383;
  assign T2383 = {4'h8/* 8*/{T138}};
  assign T2384 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2385 = T2467 && T2386;
  assign T2386 = ! T2387;
  assign T2387 = T2398 | T2388;
  assign T2388 = dramBank7_valid_received_7 & T22;
  assign T2389 = T2395 && T2390;
  assign T2390 = dramBank7_valid_received_7 || T2391;
  assign T2391 = dramBank7Port_rep_valid && T2392;
  assign T2392 = dramBank7Port_rep_tag == T2393;
  assign T2393 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign dramBank7Port_rep_tag = mainOff_dramBank7_rep_tag;
  assign mainOff_dramBank7_req_tag = dramBank7Port_req_tag;
  assign dramBank7Port_req_tag = T2394;
  assign T2394 = {6'h0/* 0*/, rThreadEncoder_io_chosen};
  assign dramBank7Port_rep_valid = mainOff_dramBank7_rep_valid;
  assign T2395 = ! T2396;
  assign T2396 = T2397 == 5'h7/* 7*/;
  assign T2397 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2398 = T2408 | T2399;
  assign T2399 = dramBank7_valid_received_6 & T73;
  assign T2400 = T2405 && T2401;
  assign T2401 = dramBank7_valid_received_6 || T2402;
  assign T2402 = dramBank7Port_rep_valid && T2403;
  assign T2403 = dramBank7Port_rep_tag == T2404;
  assign T2404 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2405 = ! T2406;
  assign T2406 = T2407 == 5'h6/* 6*/;
  assign T2407 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2408 = T2418 | T2409;
  assign T2409 = dramBank7_valid_received_5 & T84;
  assign T2410 = T2415 && T2411;
  assign T2411 = dramBank7_valid_received_5 || T2412;
  assign T2412 = dramBank7Port_rep_valid && T2413;
  assign T2413 = dramBank7Port_rep_tag == T2414;
  assign T2414 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2415 = ! T2416;
  assign T2416 = T2417 == 5'h5/* 5*/;
  assign T2417 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2418 = T2428 | T2419;
  assign T2419 = dramBank7_valid_received_4 & T95;
  assign T2420 = T2425 && T2421;
  assign T2421 = dramBank7_valid_received_4 || T2422;
  assign T2422 = dramBank7Port_rep_valid && T2423;
  assign T2423 = dramBank7Port_rep_tag == T2424;
  assign T2424 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2425 = ! T2426;
  assign T2426 = T2427 == 5'h4/* 4*/;
  assign T2427 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2428 = T2438 | T2429;
  assign T2429 = dramBank7_valid_received_3 & T106;
  assign T2430 = T2435 && T2431;
  assign T2431 = dramBank7_valid_received_3 || T2432;
  assign T2432 = dramBank7Port_rep_valid && T2433;
  assign T2433 = dramBank7Port_rep_tag == T2434;
  assign T2434 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2435 = ! T2436;
  assign T2436 = T2437 == 5'h3/* 3*/;
  assign T2437 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2438 = T2448 | T2439;
  assign T2439 = dramBank7_valid_received_2 & T117;
  assign T2440 = T2445 && T2441;
  assign T2441 = dramBank7_valid_received_2 || T2442;
  assign T2442 = dramBank7Port_rep_valid && T2443;
  assign T2443 = dramBank7Port_rep_tag == T2444;
  assign T2444 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T2445 = ! T2446;
  assign T2446 = T2447 == 5'h2/* 2*/;
  assign T2447 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2448 = T2458 | T2449;
  assign T2449 = dramBank7_valid_received_1 & T128;
  assign T2450 = T2455 && T2451;
  assign T2451 = dramBank7_valid_received_1 || T2452;
  assign T2452 = dramBank7Port_rep_valid && T2453;
  assign T2453 = dramBank7Port_rep_tag == T2454;
  assign T2454 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T2455 = ! T2456;
  assign T2456 = T2457 == 5'h1/* 1*/;
  assign T2457 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2458 = dramBank7_valid_received_0 & T138;
  assign T2459 = T2464 && T2460;
  assign T2460 = dramBank7_valid_received_0 || T2461;
  assign T2461 = dramBank7Port_rep_valid && T2462;
  assign T2462 = dramBank7Port_rep_tag == T2463;
  assign T2463 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T2464 = ! T2465;
  assign T2465 = T2466 == 5'h0/* 0*/;
  assign T2466 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2467 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T2468 = 5'h7/* 7*/ == T2469;
  assign T2469 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2470 = ! T2471;
  assign T2471 = T2472 == 5'h7/* 7*/;
  assign T2472 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2473 = T2474 || dramBank7_valid_received_7;
  assign T2474 = dramBank7Port_rep_valid && T2475;
  assign T2475 = dramBank7Port_rep_tag == T2476;
  assign T2476 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2477 = T2492 && T2478;
  assign T2478 = T2488 || T2479;
  assign T2479 = ! dramBank6PortHadValidRequest_7;
  assign T2480 = T2485 && T2481;
  assign T2481 = dramBank6PortHadValidRequest_7 || T2482;
  assign T2482 = T2483 && dramBank6Port_req_valid;
  assign T2483 = 5'h7/* 7*/ == T2484;
  assign T2484 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2485 = ! T2486;
  assign T2486 = T2487 == 5'h7/* 7*/;
  assign T2487 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2488 = T2489 || dramBank6_valid_received_7;
  assign T2489 = dramBank6Port_rep_valid && T2490;
  assign T2490 = dramBank6Port_rep_tag == T2491;
  assign T2491 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2492 = T2507 && T2493;
  assign T2493 = T2503 || T2494;
  assign T2494 = ! dramBank5PortHadValidRequest_7;
  assign T2495 = T2500 && T2496;
  assign T2496 = dramBank5PortHadValidRequest_7 || T2497;
  assign T2497 = T2498 && dramBank5Port_req_valid;
  assign T2498 = 5'h7/* 7*/ == T2499;
  assign T2499 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2500 = ! T2501;
  assign T2501 = T2502 == 5'h7/* 7*/;
  assign T2502 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2503 = T2504 || dramBank5_valid_received_7;
  assign T2504 = dramBank5Port_rep_valid && T2505;
  assign T2505 = dramBank5Port_rep_tag == T2506;
  assign T2506 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2507 = T2522 && T2508;
  assign T2508 = T2518 || T2509;
  assign T2509 = ! dramBank4PortHadValidRequest_7;
  assign T2510 = T2515 && T2511;
  assign T2511 = dramBank4PortHadValidRequest_7 || T2512;
  assign T2512 = T2513 && dramBank4Port_req_valid;
  assign T2513 = 5'h7/* 7*/ == T2514;
  assign T2514 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2515 = ! T2516;
  assign T2516 = T2517 == 5'h7/* 7*/;
  assign T2517 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2518 = T2519 || dramBank4_valid_received_7;
  assign T2519 = dramBank4Port_rep_valid && T2520;
  assign T2520 = dramBank4Port_rep_tag == T2521;
  assign T2521 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2522 = T2537 && T2523;
  assign T2523 = T2533 || T2524;
  assign T2524 = ! dramBank3PortHadValidRequest_7;
  assign T2525 = T2530 && T2526;
  assign T2526 = dramBank3PortHadValidRequest_7 || T2527;
  assign T2527 = T2528 && dramBank3Port_req_valid;
  assign T2528 = 5'h7/* 7*/ == T2529;
  assign T2529 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2530 = ! T2531;
  assign T2531 = T2532 == 5'h7/* 7*/;
  assign T2532 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2533 = T2534 || dramBank3_valid_received_7;
  assign T2534 = dramBank3Port_rep_valid && T2535;
  assign T2535 = dramBank3Port_rep_tag == T2536;
  assign T2536 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2537 = T2552 && T2538;
  assign T2538 = T2548 || T2539;
  assign T2539 = ! dramBank2PortHadValidRequest_7;
  assign T2540 = T2545 && T2541;
  assign T2541 = dramBank2PortHadValidRequest_7 || T2542;
  assign T2542 = T2543 && dramBank2Port_req_valid;
  assign T2543 = 5'h7/* 7*/ == T2544;
  assign T2544 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2545 = ! T2546;
  assign T2546 = T2547 == 5'h7/* 7*/;
  assign T2547 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2548 = T2549 || dramBank2_valid_received_7;
  assign T2549 = dramBank2Port_rep_valid && T2550;
  assign T2550 = dramBank2Port_rep_tag == T2551;
  assign T2551 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2552 = T2567 && T2553;
  assign T2553 = T2563 || T2554;
  assign T2554 = ! dramBank1PortHadValidRequest_7;
  assign T2555 = T2560 && T2556;
  assign T2556 = dramBank1PortHadValidRequest_7 || T2557;
  assign T2557 = T2558 && dramBank1Port_req_valid;
  assign T2558 = 5'h7/* 7*/ == T2559;
  assign T2559 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2560 = ! T2561;
  assign T2561 = T2562 == 5'h7/* 7*/;
  assign T2562 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2563 = T2564 || dramBank1_valid_received_7;
  assign T2564 = dramBank1Port_rep_valid && T2565;
  assign T2565 = dramBank1Port_rep_tag == T2566;
  assign T2566 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2567 = T2577 || T2568;
  assign T2568 = ! dramBank0PortHadValidRequest_7;
  assign T2569 = T2574 && T2570;
  assign T2570 = dramBank0PortHadValidRequest_7 || T2571;
  assign T2571 = T2572 && dramBank0Port_req_valid;
  assign T2572 = 5'h7/* 7*/ == T2573;
  assign T2573 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2574 = ! T2575;
  assign T2575 = T2576 == 5'h7/* 7*/;
  assign T2576 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2577 = T2578 || dramBank0_valid_received_7;
  assign T2578 = dramBank0Port_rep_valid && T2579;
  assign T2579 = dramBank0Port_rep_tag == T2580;
  assign T2580 = {5'h0/* 0*/, 5'h7/* 7*/};
  assign T2581 = subStateTh_7 == 1'h1/* 1*/;
  assign T2582 = T2702 && AllOffloadsValid_6;
  assign AllOffloadsValid_6 = T2583;
  assign T2583 = T2598 && T2584;
  assign T2584 = T2594 || T2585;
  assign T2585 = ! dramBank7PortHadValidRequest_6;
  assign T2586 = T2591 && T2587;
  assign T2587 = dramBank7PortHadValidRequest_6 || T2588;
  assign T2588 = T2589 && dramBank7Port_req_valid;
  assign T2589 = 5'h6/* 6*/ == T2590;
  assign T2590 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2591 = ! T2592;
  assign T2592 = T2593 == 5'h6/* 6*/;
  assign T2593 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2594 = T2595 || dramBank7_valid_received_6;
  assign T2595 = dramBank7Port_rep_valid && T2596;
  assign T2596 = dramBank7Port_rep_tag == T2597;
  assign T2597 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2598 = T2613 && T2599;
  assign T2599 = T2609 || T2600;
  assign T2600 = ! dramBank6PortHadValidRequest_6;
  assign T2601 = T2606 && T2602;
  assign T2602 = dramBank6PortHadValidRequest_6 || T2603;
  assign T2603 = T2604 && dramBank6Port_req_valid;
  assign T2604 = 5'h6/* 6*/ == T2605;
  assign T2605 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2606 = ! T2607;
  assign T2607 = T2608 == 5'h6/* 6*/;
  assign T2608 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2609 = T2610 || dramBank6_valid_received_6;
  assign T2610 = dramBank6Port_rep_valid && T2611;
  assign T2611 = dramBank6Port_rep_tag == T2612;
  assign T2612 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2613 = T2628 && T2614;
  assign T2614 = T2624 || T2615;
  assign T2615 = ! dramBank5PortHadValidRequest_6;
  assign T2616 = T2621 && T2617;
  assign T2617 = dramBank5PortHadValidRequest_6 || T2618;
  assign T2618 = T2619 && dramBank5Port_req_valid;
  assign T2619 = 5'h6/* 6*/ == T2620;
  assign T2620 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2621 = ! T2622;
  assign T2622 = T2623 == 5'h6/* 6*/;
  assign T2623 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2624 = T2625 || dramBank5_valid_received_6;
  assign T2625 = dramBank5Port_rep_valid && T2626;
  assign T2626 = dramBank5Port_rep_tag == T2627;
  assign T2627 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2628 = T2643 && T2629;
  assign T2629 = T2639 || T2630;
  assign T2630 = ! dramBank4PortHadValidRequest_6;
  assign T2631 = T2636 && T2632;
  assign T2632 = dramBank4PortHadValidRequest_6 || T2633;
  assign T2633 = T2634 && dramBank4Port_req_valid;
  assign T2634 = 5'h6/* 6*/ == T2635;
  assign T2635 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2636 = ! T2637;
  assign T2637 = T2638 == 5'h6/* 6*/;
  assign T2638 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2639 = T2640 || dramBank4_valid_received_6;
  assign T2640 = dramBank4Port_rep_valid && T2641;
  assign T2641 = dramBank4Port_rep_tag == T2642;
  assign T2642 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2643 = T2658 && T2644;
  assign T2644 = T2654 || T2645;
  assign T2645 = ! dramBank3PortHadValidRequest_6;
  assign T2646 = T2651 && T2647;
  assign T2647 = dramBank3PortHadValidRequest_6 || T2648;
  assign T2648 = T2649 && dramBank3Port_req_valid;
  assign T2649 = 5'h6/* 6*/ == T2650;
  assign T2650 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2651 = ! T2652;
  assign T2652 = T2653 == 5'h6/* 6*/;
  assign T2653 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2654 = T2655 || dramBank3_valid_received_6;
  assign T2655 = dramBank3Port_rep_valid && T2656;
  assign T2656 = dramBank3Port_rep_tag == T2657;
  assign T2657 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2658 = T2673 && T2659;
  assign T2659 = T2669 || T2660;
  assign T2660 = ! dramBank2PortHadValidRequest_6;
  assign T2661 = T2666 && T2662;
  assign T2662 = dramBank2PortHadValidRequest_6 || T2663;
  assign T2663 = T2664 && dramBank2Port_req_valid;
  assign T2664 = 5'h6/* 6*/ == T2665;
  assign T2665 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2666 = ! T2667;
  assign T2667 = T2668 == 5'h6/* 6*/;
  assign T2668 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2669 = T2670 || dramBank2_valid_received_6;
  assign T2670 = dramBank2Port_rep_valid && T2671;
  assign T2671 = dramBank2Port_rep_tag == T2672;
  assign T2672 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2673 = T2688 && T2674;
  assign T2674 = T2684 || T2675;
  assign T2675 = ! dramBank1PortHadValidRequest_6;
  assign T2676 = T2681 && T2677;
  assign T2677 = dramBank1PortHadValidRequest_6 || T2678;
  assign T2678 = T2679 && dramBank1Port_req_valid;
  assign T2679 = 5'h6/* 6*/ == T2680;
  assign T2680 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2681 = ! T2682;
  assign T2682 = T2683 == 5'h6/* 6*/;
  assign T2683 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2684 = T2685 || dramBank1_valid_received_6;
  assign T2685 = dramBank1Port_rep_valid && T2686;
  assign T2686 = dramBank1Port_rep_tag == T2687;
  assign T2687 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2688 = T2698 || T2689;
  assign T2689 = ! dramBank0PortHadValidRequest_6;
  assign T2690 = T2695 && T2691;
  assign T2691 = dramBank0PortHadValidRequest_6 || T2692;
  assign T2692 = T2693 && dramBank0Port_req_valid;
  assign T2693 = 5'h6/* 6*/ == T2694;
  assign T2694 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2695 = ! T2696;
  assign T2696 = T2697 == 5'h6/* 6*/;
  assign T2697 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2698 = T2699 || dramBank0_valid_received_6;
  assign T2699 = dramBank0Port_rep_valid && T2700;
  assign T2700 = dramBank0Port_rep_tag == T2701;
  assign T2701 = {5'h0/* 0*/, 5'h6/* 6*/};
  assign T2702 = subStateTh_6 == 1'h1/* 1*/;
  assign T2703 = T2823 && AllOffloadsValid_5;
  assign AllOffloadsValid_5 = T2704;
  assign T2704 = T2719 && T2705;
  assign T2705 = T2715 || T2706;
  assign T2706 = ! dramBank7PortHadValidRequest_5;
  assign T2707 = T2712 && T2708;
  assign T2708 = dramBank7PortHadValidRequest_5 || T2709;
  assign T2709 = T2710 && dramBank7Port_req_valid;
  assign T2710 = 5'h5/* 5*/ == T2711;
  assign T2711 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2712 = ! T2713;
  assign T2713 = T2714 == 5'h5/* 5*/;
  assign T2714 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2715 = T2716 || dramBank7_valid_received_5;
  assign T2716 = dramBank7Port_rep_valid && T2717;
  assign T2717 = dramBank7Port_rep_tag == T2718;
  assign T2718 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2719 = T2734 && T2720;
  assign T2720 = T2730 || T2721;
  assign T2721 = ! dramBank6PortHadValidRequest_5;
  assign T2722 = T2727 && T2723;
  assign T2723 = dramBank6PortHadValidRequest_5 || T2724;
  assign T2724 = T2725 && dramBank6Port_req_valid;
  assign T2725 = 5'h5/* 5*/ == T2726;
  assign T2726 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2727 = ! T2728;
  assign T2728 = T2729 == 5'h5/* 5*/;
  assign T2729 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2730 = T2731 || dramBank6_valid_received_5;
  assign T2731 = dramBank6Port_rep_valid && T2732;
  assign T2732 = dramBank6Port_rep_tag == T2733;
  assign T2733 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2734 = T2749 && T2735;
  assign T2735 = T2745 || T2736;
  assign T2736 = ! dramBank5PortHadValidRequest_5;
  assign T2737 = T2742 && T2738;
  assign T2738 = dramBank5PortHadValidRequest_5 || T2739;
  assign T2739 = T2740 && dramBank5Port_req_valid;
  assign T2740 = 5'h5/* 5*/ == T2741;
  assign T2741 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2742 = ! T2743;
  assign T2743 = T2744 == 5'h5/* 5*/;
  assign T2744 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2745 = T2746 || dramBank5_valid_received_5;
  assign T2746 = dramBank5Port_rep_valid && T2747;
  assign T2747 = dramBank5Port_rep_tag == T2748;
  assign T2748 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2749 = T2764 && T2750;
  assign T2750 = T2760 || T2751;
  assign T2751 = ! dramBank4PortHadValidRequest_5;
  assign T2752 = T2757 && T2753;
  assign T2753 = dramBank4PortHadValidRequest_5 || T2754;
  assign T2754 = T2755 && dramBank4Port_req_valid;
  assign T2755 = 5'h5/* 5*/ == T2756;
  assign T2756 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2757 = ! T2758;
  assign T2758 = T2759 == 5'h5/* 5*/;
  assign T2759 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2760 = T2761 || dramBank4_valid_received_5;
  assign T2761 = dramBank4Port_rep_valid && T2762;
  assign T2762 = dramBank4Port_rep_tag == T2763;
  assign T2763 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2764 = T2779 && T2765;
  assign T2765 = T2775 || T2766;
  assign T2766 = ! dramBank3PortHadValidRequest_5;
  assign T2767 = T2772 && T2768;
  assign T2768 = dramBank3PortHadValidRequest_5 || T2769;
  assign T2769 = T2770 && dramBank3Port_req_valid;
  assign T2770 = 5'h5/* 5*/ == T2771;
  assign T2771 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2772 = ! T2773;
  assign T2773 = T2774 == 5'h5/* 5*/;
  assign T2774 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2775 = T2776 || dramBank3_valid_received_5;
  assign T2776 = dramBank3Port_rep_valid && T2777;
  assign T2777 = dramBank3Port_rep_tag == T2778;
  assign T2778 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2779 = T2794 && T2780;
  assign T2780 = T2790 || T2781;
  assign T2781 = ! dramBank2PortHadValidRequest_5;
  assign T2782 = T2787 && T2783;
  assign T2783 = dramBank2PortHadValidRequest_5 || T2784;
  assign T2784 = T2785 && dramBank2Port_req_valid;
  assign T2785 = 5'h5/* 5*/ == T2786;
  assign T2786 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2787 = ! T2788;
  assign T2788 = T2789 == 5'h5/* 5*/;
  assign T2789 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2790 = T2791 || dramBank2_valid_received_5;
  assign T2791 = dramBank2Port_rep_valid && T2792;
  assign T2792 = dramBank2Port_rep_tag == T2793;
  assign T2793 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2794 = T2809 && T2795;
  assign T2795 = T2805 || T2796;
  assign T2796 = ! dramBank1PortHadValidRequest_5;
  assign T2797 = T2802 && T2798;
  assign T2798 = dramBank1PortHadValidRequest_5 || T2799;
  assign T2799 = T2800 && dramBank1Port_req_valid;
  assign T2800 = 5'h5/* 5*/ == T2801;
  assign T2801 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2802 = ! T2803;
  assign T2803 = T2804 == 5'h5/* 5*/;
  assign T2804 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2805 = T2806 || dramBank1_valid_received_5;
  assign T2806 = dramBank1Port_rep_valid && T2807;
  assign T2807 = dramBank1Port_rep_tag == T2808;
  assign T2808 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2809 = T2819 || T2810;
  assign T2810 = ! dramBank0PortHadValidRequest_5;
  assign T2811 = T2816 && T2812;
  assign T2812 = dramBank0PortHadValidRequest_5 || T2813;
  assign T2813 = T2814 && dramBank0Port_req_valid;
  assign T2814 = 5'h5/* 5*/ == T2815;
  assign T2815 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2816 = ! T2817;
  assign T2817 = T2818 == 5'h5/* 5*/;
  assign T2818 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2819 = T2820 || dramBank0_valid_received_5;
  assign T2820 = dramBank0Port_rep_valid && T2821;
  assign T2821 = dramBank0Port_rep_tag == T2822;
  assign T2822 = {5'h0/* 0*/, 5'h5/* 5*/};
  assign T2823 = subStateTh_5 == 1'h1/* 1*/;
  assign T2824 = T2944 && AllOffloadsValid_4;
  assign AllOffloadsValid_4 = T2825;
  assign T2825 = T2840 && T2826;
  assign T2826 = T2836 || T2827;
  assign T2827 = ! dramBank7PortHadValidRequest_4;
  assign T2828 = T2833 && T2829;
  assign T2829 = dramBank7PortHadValidRequest_4 || T2830;
  assign T2830 = T2831 && dramBank7Port_req_valid;
  assign T2831 = 5'h4/* 4*/ == T2832;
  assign T2832 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2833 = ! T2834;
  assign T2834 = T2835 == 5'h4/* 4*/;
  assign T2835 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2836 = T2837 || dramBank7_valid_received_4;
  assign T2837 = dramBank7Port_rep_valid && T2838;
  assign T2838 = dramBank7Port_rep_tag == T2839;
  assign T2839 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2840 = T2855 && T2841;
  assign T2841 = T2851 || T2842;
  assign T2842 = ! dramBank6PortHadValidRequest_4;
  assign T2843 = T2848 && T2844;
  assign T2844 = dramBank6PortHadValidRequest_4 || T2845;
  assign T2845 = T2846 && dramBank6Port_req_valid;
  assign T2846 = 5'h4/* 4*/ == T2847;
  assign T2847 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2848 = ! T2849;
  assign T2849 = T2850 == 5'h4/* 4*/;
  assign T2850 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2851 = T2852 || dramBank6_valid_received_4;
  assign T2852 = dramBank6Port_rep_valid && T2853;
  assign T2853 = dramBank6Port_rep_tag == T2854;
  assign T2854 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2855 = T2870 && T2856;
  assign T2856 = T2866 || T2857;
  assign T2857 = ! dramBank5PortHadValidRequest_4;
  assign T2858 = T2863 && T2859;
  assign T2859 = dramBank5PortHadValidRequest_4 || T2860;
  assign T2860 = T2861 && dramBank5Port_req_valid;
  assign T2861 = 5'h4/* 4*/ == T2862;
  assign T2862 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2863 = ! T2864;
  assign T2864 = T2865 == 5'h4/* 4*/;
  assign T2865 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2866 = T2867 || dramBank5_valid_received_4;
  assign T2867 = dramBank5Port_rep_valid && T2868;
  assign T2868 = dramBank5Port_rep_tag == T2869;
  assign T2869 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2870 = T2885 && T2871;
  assign T2871 = T2881 || T2872;
  assign T2872 = ! dramBank4PortHadValidRequest_4;
  assign T2873 = T2878 && T2874;
  assign T2874 = dramBank4PortHadValidRequest_4 || T2875;
  assign T2875 = T2876 && dramBank4Port_req_valid;
  assign T2876 = 5'h4/* 4*/ == T2877;
  assign T2877 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2878 = ! T2879;
  assign T2879 = T2880 == 5'h4/* 4*/;
  assign T2880 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2881 = T2882 || dramBank4_valid_received_4;
  assign T2882 = dramBank4Port_rep_valid && T2883;
  assign T2883 = dramBank4Port_rep_tag == T2884;
  assign T2884 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2885 = T2900 && T2886;
  assign T2886 = T2896 || T2887;
  assign T2887 = ! dramBank3PortHadValidRequest_4;
  assign T2888 = T2893 && T2889;
  assign T2889 = dramBank3PortHadValidRequest_4 || T2890;
  assign T2890 = T2891 && dramBank3Port_req_valid;
  assign T2891 = 5'h4/* 4*/ == T2892;
  assign T2892 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2893 = ! T2894;
  assign T2894 = T2895 == 5'h4/* 4*/;
  assign T2895 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2896 = T2897 || dramBank3_valid_received_4;
  assign T2897 = dramBank3Port_rep_valid && T2898;
  assign T2898 = dramBank3Port_rep_tag == T2899;
  assign T2899 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2900 = T2915 && T2901;
  assign T2901 = T2911 || T2902;
  assign T2902 = ! dramBank2PortHadValidRequest_4;
  assign T2903 = T2908 && T2904;
  assign T2904 = dramBank2PortHadValidRequest_4 || T2905;
  assign T2905 = T2906 && dramBank2Port_req_valid;
  assign T2906 = 5'h4/* 4*/ == T2907;
  assign T2907 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2908 = ! T2909;
  assign T2909 = T2910 == 5'h4/* 4*/;
  assign T2910 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2911 = T2912 || dramBank2_valid_received_4;
  assign T2912 = dramBank2Port_rep_valid && T2913;
  assign T2913 = dramBank2Port_rep_tag == T2914;
  assign T2914 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2915 = T2930 && T2916;
  assign T2916 = T2926 || T2917;
  assign T2917 = ! dramBank1PortHadValidRequest_4;
  assign T2918 = T2923 && T2919;
  assign T2919 = dramBank1PortHadValidRequest_4 || T2920;
  assign T2920 = T2921 && dramBank1Port_req_valid;
  assign T2921 = 5'h4/* 4*/ == T2922;
  assign T2922 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2923 = ! T2924;
  assign T2924 = T2925 == 5'h4/* 4*/;
  assign T2925 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2926 = T2927 || dramBank1_valid_received_4;
  assign T2927 = dramBank1Port_rep_valid && T2928;
  assign T2928 = dramBank1Port_rep_tag == T2929;
  assign T2929 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2930 = T2940 || T2931;
  assign T2931 = ! dramBank0PortHadValidRequest_4;
  assign T2932 = T2937 && T2933;
  assign T2933 = dramBank0PortHadValidRequest_4 || T2934;
  assign T2934 = T2935 && dramBank0Port_req_valid;
  assign T2935 = 5'h4/* 4*/ == T2936;
  assign T2936 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2937 = ! T2938;
  assign T2938 = T2939 == 5'h4/* 4*/;
  assign T2939 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2940 = T2941 || dramBank0_valid_received_4;
  assign T2941 = dramBank0Port_rep_valid && T2942;
  assign T2942 = dramBank0Port_rep_tag == T2943;
  assign T2943 = {5'h0/* 0*/, 5'h4/* 4*/};
  assign T2944 = subStateTh_4 == 1'h1/* 1*/;
  assign T2945 = T3065 && AllOffloadsValid_3;
  assign AllOffloadsValid_3 = T2946;
  assign T2946 = T2961 && T2947;
  assign T2947 = T2957 || T2948;
  assign T2948 = ! dramBank7PortHadValidRequest_3;
  assign T2949 = T2954 && T2950;
  assign T2950 = dramBank7PortHadValidRequest_3 || T2951;
  assign T2951 = T2952 && dramBank7Port_req_valid;
  assign T2952 = 5'h3/* 3*/ == T2953;
  assign T2953 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2954 = ! T2955;
  assign T2955 = T2956 == 5'h3/* 3*/;
  assign T2956 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2957 = T2958 || dramBank7_valid_received_3;
  assign T2958 = dramBank7Port_rep_valid && T2959;
  assign T2959 = dramBank7Port_rep_tag == T2960;
  assign T2960 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2961 = T2976 && T2962;
  assign T2962 = T2972 || T2963;
  assign T2963 = ! dramBank6PortHadValidRequest_3;
  assign T2964 = T2969 && T2965;
  assign T2965 = dramBank6PortHadValidRequest_3 || T2966;
  assign T2966 = T2967 && dramBank6Port_req_valid;
  assign T2967 = 5'h3/* 3*/ == T2968;
  assign T2968 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2969 = ! T2970;
  assign T2970 = T2971 == 5'h3/* 3*/;
  assign T2971 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2972 = T2973 || dramBank6_valid_received_3;
  assign T2973 = dramBank6Port_rep_valid && T2974;
  assign T2974 = dramBank6Port_rep_tag == T2975;
  assign T2975 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2976 = T2991 && T2977;
  assign T2977 = T2987 || T2978;
  assign T2978 = ! dramBank5PortHadValidRequest_3;
  assign T2979 = T2984 && T2980;
  assign T2980 = dramBank5PortHadValidRequest_3 || T2981;
  assign T2981 = T2982 && dramBank5Port_req_valid;
  assign T2982 = 5'h3/* 3*/ == T2983;
  assign T2983 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2984 = ! T2985;
  assign T2985 = T2986 == 5'h3/* 3*/;
  assign T2986 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T2987 = T2988 || dramBank5_valid_received_3;
  assign T2988 = dramBank5Port_rep_valid && T2989;
  assign T2989 = dramBank5Port_rep_tag == T2990;
  assign T2990 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T2991 = T3006 && T2992;
  assign T2992 = T3002 || T2993;
  assign T2993 = ! dramBank4PortHadValidRequest_3;
  assign T2994 = T2999 && T2995;
  assign T2995 = dramBank4PortHadValidRequest_3 || T2996;
  assign T2996 = T2997 && dramBank4Port_req_valid;
  assign T2997 = 5'h3/* 3*/ == T2998;
  assign T2998 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T2999 = ! T3000;
  assign T3000 = T3001 == 5'h3/* 3*/;
  assign T3001 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3002 = T3003 || dramBank4_valid_received_3;
  assign T3003 = dramBank4Port_rep_valid && T3004;
  assign T3004 = dramBank4Port_rep_tag == T3005;
  assign T3005 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3006 = T3021 && T3007;
  assign T3007 = T3017 || T3008;
  assign T3008 = ! dramBank3PortHadValidRequest_3;
  assign T3009 = T3014 && T3010;
  assign T3010 = dramBank3PortHadValidRequest_3 || T3011;
  assign T3011 = T3012 && dramBank3Port_req_valid;
  assign T3012 = 5'h3/* 3*/ == T3013;
  assign T3013 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3014 = ! T3015;
  assign T3015 = T3016 == 5'h3/* 3*/;
  assign T3016 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3017 = T3018 || dramBank3_valid_received_3;
  assign T3018 = dramBank3Port_rep_valid && T3019;
  assign T3019 = dramBank3Port_rep_tag == T3020;
  assign T3020 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3021 = T3036 && T3022;
  assign T3022 = T3032 || T3023;
  assign T3023 = ! dramBank2PortHadValidRequest_3;
  assign T3024 = T3029 && T3025;
  assign T3025 = dramBank2PortHadValidRequest_3 || T3026;
  assign T3026 = T3027 && dramBank2Port_req_valid;
  assign T3027 = 5'h3/* 3*/ == T3028;
  assign T3028 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3029 = ! T3030;
  assign T3030 = T3031 == 5'h3/* 3*/;
  assign T3031 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3032 = T3033 || dramBank2_valid_received_3;
  assign T3033 = dramBank2Port_rep_valid && T3034;
  assign T3034 = dramBank2Port_rep_tag == T3035;
  assign T3035 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3036 = T3051 && T3037;
  assign T3037 = T3047 || T3038;
  assign T3038 = ! dramBank1PortHadValidRequest_3;
  assign T3039 = T3044 && T3040;
  assign T3040 = dramBank1PortHadValidRequest_3 || T3041;
  assign T3041 = T3042 && dramBank1Port_req_valid;
  assign T3042 = 5'h3/* 3*/ == T3043;
  assign T3043 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3044 = ! T3045;
  assign T3045 = T3046 == 5'h3/* 3*/;
  assign T3046 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3047 = T3048 || dramBank1_valid_received_3;
  assign T3048 = dramBank1Port_rep_valid && T3049;
  assign T3049 = dramBank1Port_rep_tag == T3050;
  assign T3050 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3051 = T3061 || T3052;
  assign T3052 = ! dramBank0PortHadValidRequest_3;
  assign T3053 = T3058 && T3054;
  assign T3054 = dramBank0PortHadValidRequest_3 || T3055;
  assign T3055 = T3056 && dramBank0Port_req_valid;
  assign T3056 = 5'h3/* 3*/ == T3057;
  assign T3057 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3058 = ! T3059;
  assign T3059 = T3060 == 5'h3/* 3*/;
  assign T3060 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3061 = T3062 || dramBank0_valid_received_3;
  assign T3062 = dramBank0Port_rep_valid && T3063;
  assign T3063 = dramBank0Port_rep_tag == T3064;
  assign T3064 = {5'h0/* 0*/, 5'h3/* 3*/};
  assign T3065 = subStateTh_3 == 1'h1/* 1*/;
  assign T3066 = T3186 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T3067;
  assign T3067 = T3082 && T3068;
  assign T3068 = T3078 || T3069;
  assign T3069 = ! dramBank7PortHadValidRequest_2;
  assign T3070 = T3075 && T3071;
  assign T3071 = dramBank7PortHadValidRequest_2 || T3072;
  assign T3072 = T3073 && dramBank7Port_req_valid;
  assign T3073 = 5'h2/* 2*/ == T3074;
  assign T3074 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3075 = ! T3076;
  assign T3076 = T3077 == 5'h2/* 2*/;
  assign T3077 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3078 = T3079 || dramBank7_valid_received_2;
  assign T3079 = dramBank7Port_rep_valid && T3080;
  assign T3080 = dramBank7Port_rep_tag == T3081;
  assign T3081 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3082 = T3097 && T3083;
  assign T3083 = T3093 || T3084;
  assign T3084 = ! dramBank6PortHadValidRequest_2;
  assign T3085 = T3090 && T3086;
  assign T3086 = dramBank6PortHadValidRequest_2 || T3087;
  assign T3087 = T3088 && dramBank6Port_req_valid;
  assign T3088 = 5'h2/* 2*/ == T3089;
  assign T3089 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3090 = ! T3091;
  assign T3091 = T3092 == 5'h2/* 2*/;
  assign T3092 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3093 = T3094 || dramBank6_valid_received_2;
  assign T3094 = dramBank6Port_rep_valid && T3095;
  assign T3095 = dramBank6Port_rep_tag == T3096;
  assign T3096 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3097 = T3112 && T3098;
  assign T3098 = T3108 || T3099;
  assign T3099 = ! dramBank5PortHadValidRequest_2;
  assign T3100 = T3105 && T3101;
  assign T3101 = dramBank5PortHadValidRequest_2 || T3102;
  assign T3102 = T3103 && dramBank5Port_req_valid;
  assign T3103 = 5'h2/* 2*/ == T3104;
  assign T3104 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3105 = ! T3106;
  assign T3106 = T3107 == 5'h2/* 2*/;
  assign T3107 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3108 = T3109 || dramBank5_valid_received_2;
  assign T3109 = dramBank5Port_rep_valid && T3110;
  assign T3110 = dramBank5Port_rep_tag == T3111;
  assign T3111 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3112 = T3127 && T3113;
  assign T3113 = T3123 || T3114;
  assign T3114 = ! dramBank4PortHadValidRequest_2;
  assign T3115 = T3120 && T3116;
  assign T3116 = dramBank4PortHadValidRequest_2 || T3117;
  assign T3117 = T3118 && dramBank4Port_req_valid;
  assign T3118 = 5'h2/* 2*/ == T3119;
  assign T3119 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3120 = ! T3121;
  assign T3121 = T3122 == 5'h2/* 2*/;
  assign T3122 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3123 = T3124 || dramBank4_valid_received_2;
  assign T3124 = dramBank4Port_rep_valid && T3125;
  assign T3125 = dramBank4Port_rep_tag == T3126;
  assign T3126 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3127 = T3142 && T3128;
  assign T3128 = T3138 || T3129;
  assign T3129 = ! dramBank3PortHadValidRequest_2;
  assign T3130 = T3135 && T3131;
  assign T3131 = dramBank3PortHadValidRequest_2 || T3132;
  assign T3132 = T3133 && dramBank3Port_req_valid;
  assign T3133 = 5'h2/* 2*/ == T3134;
  assign T3134 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3135 = ! T3136;
  assign T3136 = T3137 == 5'h2/* 2*/;
  assign T3137 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3138 = T3139 || dramBank3_valid_received_2;
  assign T3139 = dramBank3Port_rep_valid && T3140;
  assign T3140 = dramBank3Port_rep_tag == T3141;
  assign T3141 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3142 = T3157 && T3143;
  assign T3143 = T3153 || T3144;
  assign T3144 = ! dramBank2PortHadValidRequest_2;
  assign T3145 = T3150 && T3146;
  assign T3146 = dramBank2PortHadValidRequest_2 || T3147;
  assign T3147 = T3148 && dramBank2Port_req_valid;
  assign T3148 = 5'h2/* 2*/ == T3149;
  assign T3149 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3150 = ! T3151;
  assign T3151 = T3152 == 5'h2/* 2*/;
  assign T3152 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3153 = T3154 || dramBank2_valid_received_2;
  assign T3154 = dramBank2Port_rep_valid && T3155;
  assign T3155 = dramBank2Port_rep_tag == T3156;
  assign T3156 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3157 = T3172 && T3158;
  assign T3158 = T3168 || T3159;
  assign T3159 = ! dramBank1PortHadValidRequest_2;
  assign T3160 = T3165 && T3161;
  assign T3161 = dramBank1PortHadValidRequest_2 || T3162;
  assign T3162 = T3163 && dramBank1Port_req_valid;
  assign T3163 = 5'h2/* 2*/ == T3164;
  assign T3164 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3165 = ! T3166;
  assign T3166 = T3167 == 5'h2/* 2*/;
  assign T3167 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3168 = T3169 || dramBank1_valid_received_2;
  assign T3169 = dramBank1Port_rep_valid && T3170;
  assign T3170 = dramBank1Port_rep_tag == T3171;
  assign T3171 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3172 = T3182 || T3173;
  assign T3173 = ! dramBank0PortHadValidRequest_2;
  assign T3174 = T3179 && T3175;
  assign T3175 = dramBank0PortHadValidRequest_2 || T3176;
  assign T3176 = T3177 && dramBank0Port_req_valid;
  assign T3177 = 5'h2/* 2*/ == T3178;
  assign T3178 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3179 = ! T3180;
  assign T3180 = T3181 == 5'h2/* 2*/;
  assign T3181 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3182 = T3183 || dramBank0_valid_received_2;
  assign T3183 = dramBank0Port_rep_valid && T3184;
  assign T3184 = dramBank0Port_rep_tag == T3185;
  assign T3185 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T3186 = subStateTh_2 == 1'h1/* 1*/;
  assign T3187 = T3307 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T3188;
  assign T3188 = T3203 && T3189;
  assign T3189 = T3199 || T3190;
  assign T3190 = ! dramBank7PortHadValidRequest_1;
  assign T3191 = T3196 && T3192;
  assign T3192 = dramBank7PortHadValidRequest_1 || T3193;
  assign T3193 = T3194 && dramBank7Port_req_valid;
  assign T3194 = 5'h1/* 1*/ == T3195;
  assign T3195 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3196 = ! T3197;
  assign T3197 = T3198 == 5'h1/* 1*/;
  assign T3198 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3199 = T3200 || dramBank7_valid_received_1;
  assign T3200 = dramBank7Port_rep_valid && T3201;
  assign T3201 = dramBank7Port_rep_tag == T3202;
  assign T3202 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3203 = T3218 && T3204;
  assign T3204 = T3214 || T3205;
  assign T3205 = ! dramBank6PortHadValidRequest_1;
  assign T3206 = T3211 && T3207;
  assign T3207 = dramBank6PortHadValidRequest_1 || T3208;
  assign T3208 = T3209 && dramBank6Port_req_valid;
  assign T3209 = 5'h1/* 1*/ == T3210;
  assign T3210 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3211 = ! T3212;
  assign T3212 = T3213 == 5'h1/* 1*/;
  assign T3213 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3214 = T3215 || dramBank6_valid_received_1;
  assign T3215 = dramBank6Port_rep_valid && T3216;
  assign T3216 = dramBank6Port_rep_tag == T3217;
  assign T3217 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3218 = T3233 && T3219;
  assign T3219 = T3229 || T3220;
  assign T3220 = ! dramBank5PortHadValidRequest_1;
  assign T3221 = T3226 && T3222;
  assign T3222 = dramBank5PortHadValidRequest_1 || T3223;
  assign T3223 = T3224 && dramBank5Port_req_valid;
  assign T3224 = 5'h1/* 1*/ == T3225;
  assign T3225 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3226 = ! T3227;
  assign T3227 = T3228 == 5'h1/* 1*/;
  assign T3228 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3229 = T3230 || dramBank5_valid_received_1;
  assign T3230 = dramBank5Port_rep_valid && T3231;
  assign T3231 = dramBank5Port_rep_tag == T3232;
  assign T3232 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3233 = T3248 && T3234;
  assign T3234 = T3244 || T3235;
  assign T3235 = ! dramBank4PortHadValidRequest_1;
  assign T3236 = T3241 && T3237;
  assign T3237 = dramBank4PortHadValidRequest_1 || T3238;
  assign T3238 = T3239 && dramBank4Port_req_valid;
  assign T3239 = 5'h1/* 1*/ == T3240;
  assign T3240 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3241 = ! T3242;
  assign T3242 = T3243 == 5'h1/* 1*/;
  assign T3243 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3244 = T3245 || dramBank4_valid_received_1;
  assign T3245 = dramBank4Port_rep_valid && T3246;
  assign T3246 = dramBank4Port_rep_tag == T3247;
  assign T3247 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3248 = T3263 && T3249;
  assign T3249 = T3259 || T3250;
  assign T3250 = ! dramBank3PortHadValidRequest_1;
  assign T3251 = T3256 && T3252;
  assign T3252 = dramBank3PortHadValidRequest_1 || T3253;
  assign T3253 = T3254 && dramBank3Port_req_valid;
  assign T3254 = 5'h1/* 1*/ == T3255;
  assign T3255 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3256 = ! T3257;
  assign T3257 = T3258 == 5'h1/* 1*/;
  assign T3258 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3259 = T3260 || dramBank3_valid_received_1;
  assign T3260 = dramBank3Port_rep_valid && T3261;
  assign T3261 = dramBank3Port_rep_tag == T3262;
  assign T3262 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3263 = T3278 && T3264;
  assign T3264 = T3274 || T3265;
  assign T3265 = ! dramBank2PortHadValidRequest_1;
  assign T3266 = T3271 && T3267;
  assign T3267 = dramBank2PortHadValidRequest_1 || T3268;
  assign T3268 = T3269 && dramBank2Port_req_valid;
  assign T3269 = 5'h1/* 1*/ == T3270;
  assign T3270 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3271 = ! T3272;
  assign T3272 = T3273 == 5'h1/* 1*/;
  assign T3273 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3274 = T3275 || dramBank2_valid_received_1;
  assign T3275 = dramBank2Port_rep_valid && T3276;
  assign T3276 = dramBank2Port_rep_tag == T3277;
  assign T3277 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3278 = T3293 && T3279;
  assign T3279 = T3289 || T3280;
  assign T3280 = ! dramBank1PortHadValidRequest_1;
  assign T3281 = T3286 && T3282;
  assign T3282 = dramBank1PortHadValidRequest_1 || T3283;
  assign T3283 = T3284 && dramBank1Port_req_valid;
  assign T3284 = 5'h1/* 1*/ == T3285;
  assign T3285 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3286 = ! T3287;
  assign T3287 = T3288 == 5'h1/* 1*/;
  assign T3288 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3289 = T3290 || dramBank1_valid_received_1;
  assign T3290 = dramBank1Port_rep_valid && T3291;
  assign T3291 = dramBank1Port_rep_tag == T3292;
  assign T3292 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3293 = T3303 || T3294;
  assign T3294 = ! dramBank0PortHadValidRequest_1;
  assign T3295 = T3300 && T3296;
  assign T3296 = dramBank0PortHadValidRequest_1 || T3297;
  assign T3297 = T3298 && dramBank0Port_req_valid;
  assign T3298 = 5'h1/* 1*/ == T3299;
  assign T3299 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3300 = ! T3301;
  assign T3301 = T3302 == 5'h1/* 1*/;
  assign T3302 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3303 = T3304 || dramBank0_valid_received_1;
  assign T3304 = dramBank0Port_rep_valid && T3305;
  assign T3305 = dramBank0Port_rep_tag == T3306;
  assign T3306 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T3307 = subStateTh_1 == 1'h1/* 1*/;
  assign T3308 = T3428 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T3309;
  assign T3309 = T3324 && T3310;
  assign T3310 = T3320 || T3311;
  assign T3311 = ! dramBank7PortHadValidRequest_0;
  assign T3312 = T3317 && T3313;
  assign T3313 = dramBank7PortHadValidRequest_0 || T3314;
  assign T3314 = T3315 && dramBank7Port_req_valid;
  assign T3315 = 5'h0/* 0*/ == T3316;
  assign T3316 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3317 = ! T3318;
  assign T3318 = T3319 == 5'h0/* 0*/;
  assign T3319 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3320 = T3321 || dramBank7_valid_received_0;
  assign T3321 = dramBank7Port_rep_valid && T3322;
  assign T3322 = dramBank7Port_rep_tag == T3323;
  assign T3323 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3324 = T3339 && T3325;
  assign T3325 = T3335 || T3326;
  assign T3326 = ! dramBank6PortHadValidRequest_0;
  assign T3327 = T3332 && T3328;
  assign T3328 = dramBank6PortHadValidRequest_0 || T3329;
  assign T3329 = T3330 && dramBank6Port_req_valid;
  assign T3330 = 5'h0/* 0*/ == T3331;
  assign T3331 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3332 = ! T3333;
  assign T3333 = T3334 == 5'h0/* 0*/;
  assign T3334 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3335 = T3336 || dramBank6_valid_received_0;
  assign T3336 = dramBank6Port_rep_valid && T3337;
  assign T3337 = dramBank6Port_rep_tag == T3338;
  assign T3338 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3339 = T3354 && T3340;
  assign T3340 = T3350 || T3341;
  assign T3341 = ! dramBank5PortHadValidRequest_0;
  assign T3342 = T3347 && T3343;
  assign T3343 = dramBank5PortHadValidRequest_0 || T3344;
  assign T3344 = T3345 && dramBank5Port_req_valid;
  assign T3345 = 5'h0/* 0*/ == T3346;
  assign T3346 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3347 = ! T3348;
  assign T3348 = T3349 == 5'h0/* 0*/;
  assign T3349 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3350 = T3351 || dramBank5_valid_received_0;
  assign T3351 = dramBank5Port_rep_valid && T3352;
  assign T3352 = dramBank5Port_rep_tag == T3353;
  assign T3353 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3354 = T3369 && T3355;
  assign T3355 = T3365 || T3356;
  assign T3356 = ! dramBank4PortHadValidRequest_0;
  assign T3357 = T3362 && T3358;
  assign T3358 = dramBank4PortHadValidRequest_0 || T3359;
  assign T3359 = T3360 && dramBank4Port_req_valid;
  assign T3360 = 5'h0/* 0*/ == T3361;
  assign T3361 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3362 = ! T3363;
  assign T3363 = T3364 == 5'h0/* 0*/;
  assign T3364 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3365 = T3366 || dramBank4_valid_received_0;
  assign T3366 = dramBank4Port_rep_valid && T3367;
  assign T3367 = dramBank4Port_rep_tag == T3368;
  assign T3368 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3369 = T3384 && T3370;
  assign T3370 = T3380 || T3371;
  assign T3371 = ! dramBank3PortHadValidRequest_0;
  assign T3372 = T3377 && T3373;
  assign T3373 = dramBank3PortHadValidRequest_0 || T3374;
  assign T3374 = T3375 && dramBank3Port_req_valid;
  assign T3375 = 5'h0/* 0*/ == T3376;
  assign T3376 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3377 = ! T3378;
  assign T3378 = T3379 == 5'h0/* 0*/;
  assign T3379 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3380 = T3381 || dramBank3_valid_received_0;
  assign T3381 = dramBank3Port_rep_valid && T3382;
  assign T3382 = dramBank3Port_rep_tag == T3383;
  assign T3383 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3384 = T3399 && T3385;
  assign T3385 = T3395 || T3386;
  assign T3386 = ! dramBank2PortHadValidRequest_0;
  assign T3387 = T3392 && T3388;
  assign T3388 = dramBank2PortHadValidRequest_0 || T3389;
  assign T3389 = T3390 && dramBank2Port_req_valid;
  assign T3390 = 5'h0/* 0*/ == T3391;
  assign T3391 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3392 = ! T3393;
  assign T3393 = T3394 == 5'h0/* 0*/;
  assign T3394 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3395 = T3396 || dramBank2_valid_received_0;
  assign T3396 = dramBank2Port_rep_valid && T3397;
  assign T3397 = dramBank2Port_rep_tag == T3398;
  assign T3398 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3399 = T3414 && T3400;
  assign T3400 = T3410 || T3401;
  assign T3401 = ! dramBank1PortHadValidRequest_0;
  assign T3402 = T3407 && T3403;
  assign T3403 = dramBank1PortHadValidRequest_0 || T3404;
  assign T3404 = T3405 && dramBank1Port_req_valid;
  assign T3405 = 5'h0/* 0*/ == T3406;
  assign T3406 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3407 = ! T3408;
  assign T3408 = T3409 == 5'h0/* 0*/;
  assign T3409 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3410 = T3411 || dramBank1_valid_received_0;
  assign T3411 = dramBank1Port_rep_valid && T3412;
  assign T3412 = dramBank1Port_rep_tag == T3413;
  assign T3413 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3414 = T3424 || T3415;
  assign T3415 = ! dramBank0PortHadValidRequest_0;
  assign T3416 = T3421 && T3417;
  assign T3417 = dramBank0PortHadValidRequest_0 || T3418;
  assign T3418 = T3419 && dramBank0Port_req_valid;
  assign T3419 = 5'h0/* 0*/ == T3420;
  assign T3420 = {1'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T3421 = ! T3422;
  assign T3422 = T3423 == 5'h0/* 0*/;
  assign T3423 = {1'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T3424 = T3425 || dramBank0_valid_received_0;
  assign T3425 = dramBank0Port_rep_valid && T3426;
  assign T3426 = dramBank0Port_rep_tag == T3427;
  assign T3427 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T3428 = subStateTh_0 == 1'h1/* 1*/;
  assign T3429 = vThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign T3430 = T3431 || T1534;
  assign T3431 = T3432 || T1536;
  assign T3432 = T3433 || T1538;
  assign T3433 = T3434 || T1540;
  assign T3434 = T3435 || T1542;
  assign T3435 = T3436 || T1544;
  assign T3436 = T3437 || T1546;
  assign T3437 = T3438 || T1547;
  assign T3438 = T3440 || T3439;
  assign T3439 = T830 && T5;
  assign T3440 = T3441 || T936;
  assign T3441 = T3443 || T3442;
  assign T3442 = T997 && T5;
  assign T3443 = T3444 || T1008;
  assign T3444 = T3446 || T3445;
  assign T3445 = T1069 && T5;
  assign T3446 = T3447 || T1080;
  assign T3447 = T3449 || T3448;
  assign T3448 = T1141 && T5;
  assign T3449 = T3450 || T1152;
  assign T3450 = T3452 || T3451;
  assign T3451 = T1213 && T5;
  assign T3452 = T3453 || T1224;
  assign T3453 = T3455 || T3454;
  assign T3454 = T1285 && T5;
  assign T3455 = T3456 || T1296;
  assign T3456 = T3458 || T3457;
  assign T3457 = T1357 && T5;
  assign T3458 = T3459 || T1368;
  assign T3459 = T3461 || T3460;
  assign T3460 = T1429 && T5;
  assign T3461 = T3462 || T1440;
  assign T3462 = T3464 || T3463;
  assign T3463 = T1501 && T5;
  assign T3464 = T839 || T3465;
  assign T3465 = T1504 && T22;
  assign T3466 = T3504 ? 8'hff/* 255*/ : T3467;
  assign T3467 = T3439 ? T3503 : T3468;
  assign T3468 = T936 ? T3502 : T3469;
  assign T3469 = T3442 ? T3501 : T3470;
  assign T3470 = T1008 ? T3500 : T3471;
  assign T3471 = T3445 ? T3499 : T3472;
  assign T3472 = T1080 ? T3498 : T3473;
  assign T3473 = T3448 ? T3497 : T3474;
  assign T3474 = T1152 ? T3496 : T3475;
  assign T3475 = T3451 ? T3495 : T3476;
  assign T3476 = T1224 ? T3494 : T3477;
  assign T3477 = T3454 ? T3493 : T3478;
  assign T3478 = T1296 ? T3492 : T3479;
  assign T3479 = T3457 ? T3491 : T3480;
  assign T3480 = T1368 ? T3490 : T3481;
  assign T3481 = T3460 ? T3489 : T3482;
  assign T3482 = T1440 ? T3488 : T3483;
  assign T3483 = T3463 ? T3487 : T3484;
  assign T3484 = T3465 ? T1529 : T3485;
  assign T3485 = T839 ? T3486 : State_7;
  assign T3486 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T3487 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3488 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T3489 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3490 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T3491 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3492 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T3493 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T3495 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3496 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T3497 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3498 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T3499 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3500 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T3501 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3502 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T3503 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T3504 = T3505 || T4;
  assign T3505 = T3506 || T1534;
  assign T3506 = T3507 || T1536;
  assign T3507 = T3508 || T1538;
  assign T3508 = T3509 || T1540;
  assign T3509 = T3510 || T1542;
  assign T3510 = T3511 || T1544;
  assign T3511 = T1547 || T1546;
  assign T3512 = subStateTh_7 == 1'h0/* 0*/;
  assign T3513 = T3515 && T3514;
  assign T3514 = State_6 == 8'h0/* 0*/;
  assign T3515 = subStateTh_6 == 1'h0/* 0*/;
  assign T3516 = T3518 && T3517;
  assign T3517 = State_5 == 8'h0/* 0*/;
  assign T3518 = subStateTh_5 == 1'h0/* 0*/;
  assign T3519 = T3521 && T3520;
  assign T3520 = State_4 == 8'h0/* 0*/;
  assign T3521 = subStateTh_4 == 1'h0/* 0*/;
  assign T3522 = T3524 && T3523;
  assign T3523 = State_3 == 8'h0/* 0*/;
  assign T3524 = subStateTh_3 == 1'h0/* 0*/;
  assign T3525 = T3527 && T3526;
  assign T3526 = State_2 == 8'h0/* 0*/;
  assign T3527 = subStateTh_2 == 1'h0/* 0*/;
  assign T3528 = T3530 && T3529;
  assign T3529 = State_1 == 8'h0/* 0*/;
  assign T3530 = subStateTh_1 == 1'h0/* 0*/;
  assign T3531 = T3533 && T3532;
  assign T3532 = State_0 == 8'h0/* 0*/;
  assign T3533 = subStateTh_0 == 1'h0/* 0*/;
  assign T3534 = sThreadEncoder_io_chosen != 4'h8/* 8*/;
  assign io_out_tag = T3535;
  assign T3535 = T3539 | T3536;
  assign T3536 = inputTag_7 & T3537;
  assign T3537 = {4'ha/* 10*/{T22}};
  assign T3538 = T839 ? io_in_tag : inputTag_7;
  assign T3539 = T3543 | T3540;
  assign T3540 = inputTag_6 & T3541;
  assign T3541 = {4'ha/* 10*/{T73}};
  assign T3542 = T849 ? io_in_tag : inputTag_6;
  assign T3543 = T3547 | T3544;
  assign T3544 = inputTag_5 & T3545;
  assign T3545 = {4'ha/* 10*/{T84}};
  assign T3546 = T855 ? io_in_tag : inputTag_5;
  assign T3547 = T3551 | T3548;
  assign T3548 = inputTag_4 & T3549;
  assign T3549 = {4'ha/* 10*/{T95}};
  assign T3550 = T862 ? io_in_tag : inputTag_4;
  assign T3551 = T3555 | T3552;
  assign T3552 = inputTag_3 & T3553;
  assign T3553 = {4'ha/* 10*/{T106}};
  assign T3554 = T869 ? io_in_tag : inputTag_3;
  assign T3555 = T3559 | T3556;
  assign T3556 = inputTag_2 & T3557;
  assign T3557 = {4'ha/* 10*/{T117}};
  assign T3558 = T876 ? io_in_tag : inputTag_2;
  assign T3559 = T3563 | T3560;
  assign T3560 = inputTag_1 & T3561;
  assign T3561 = {4'ha/* 10*/{T128}};
  assign T3562 = T883 ? io_in_tag : inputTag_1;
  assign T3563 = inputTag_0 & T3564;
  assign T3564 = {4'ha/* 10*/{T138}};
  assign T3565 = T889 ? io_in_tag : inputTag_0;
  assign io_out_valid = T3566;
  assign T3566 = T3568 && T3567;
  assign T3567 = T19 == 8'hff/* 255*/;
  assign T3568 = rThreadEncoder_io_chosen != 4'h8/* 8*/;
  RREncode_59 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T2351 ),
       .io_valid_1( T2339 ),
       .io_valid_2( T2327 ),
       .io_valid_3( T2315 ),
       .io_valid_4( T2303 ),
       .io_valid_5( T2291 ),
       .io_valid_6( T755 ),
       .io_valid_7( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T2363 ));
  RREncode_60 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T3308 ),
       .io_valid_1( T3187 ),
       .io_valid_2( T3066 ),
       .io_valid_3( T2945 ),
       .io_valid_4( T2824 ),
       .io_valid_5( T2703 ),
       .io_valid_6( T2582 ),
       .io_valid_7( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T3429 ));
  RREncode_61 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T3531 ),
       .io_valid_1( T3528 ),
       .io_valid_2( T3525 ),
       .io_valid_3( T3522 ),
       .io_valid_4( T3519 ),
       .io_valid_5( T3516 ),
       .io_valid_6( T3513 ),
       .io_valid_7( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T3534 ));

  always @(posedge clk) begin
    if(reset) begin
      State_7 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_7 <= T3466;
    end
    dramBank7PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_7 <= reset ? 1'h0/* 0*/ : T26;
    dramBank7PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T42;
    dramBank7_ready_received <= reset ? 1'h0/* 0*/ : T46;
    dramBank6_valid_received_7 <= reset ? 1'h0/* 0*/ : T62;
    dramBank6_valid_received_6 <= reset ? 1'h0/* 0*/ : T74;
    dramBank6_valid_received_5 <= reset ? 1'h0/* 0*/ : T85;
    dramBank6_valid_received_4 <= reset ? 1'h0/* 0*/ : T96;
    dramBank6_valid_received_3 <= reset ? 1'h0/* 0*/ : T107;
    dramBank6_valid_received_2 <= reset ? 1'h0/* 0*/ : T118;
    dramBank6_valid_received_1 <= reset ? 1'h0/* 0*/ : T129;
    dramBank6_valid_received_0 <= reset ? 1'h0/* 0*/ : T139;
    dramBank6PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T149;
    dramBank6_ready_received <= reset ? 1'h0/* 0*/ : T153;
    dramBank5_valid_received_7 <= reset ? 1'h0/* 0*/ : T169;
    dramBank5_valid_received_6 <= reset ? 1'h0/* 0*/ : T180;
    dramBank5_valid_received_5 <= reset ? 1'h0/* 0*/ : T190;
    dramBank5_valid_received_4 <= reset ? 1'h0/* 0*/ : T200;
    dramBank5_valid_received_3 <= reset ? 1'h0/* 0*/ : T210;
    dramBank5_valid_received_2 <= reset ? 1'h0/* 0*/ : T220;
    dramBank5_valid_received_1 <= reset ? 1'h0/* 0*/ : T230;
    dramBank5_valid_received_0 <= reset ? 1'h0/* 0*/ : T239;
    dramBank5PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T249;
    dramBank5_ready_received <= reset ? 1'h0/* 0*/ : T253;
    dramBank4_valid_received_7 <= reset ? 1'h0/* 0*/ : T269;
    dramBank4_valid_received_6 <= reset ? 1'h0/* 0*/ : T280;
    dramBank4_valid_received_5 <= reset ? 1'h0/* 0*/ : T290;
    dramBank4_valid_received_4 <= reset ? 1'h0/* 0*/ : T300;
    dramBank4_valid_received_3 <= reset ? 1'h0/* 0*/ : T310;
    dramBank4_valid_received_2 <= reset ? 1'h0/* 0*/ : T320;
    dramBank4_valid_received_1 <= reset ? 1'h0/* 0*/ : T330;
    dramBank4_valid_received_0 <= reset ? 1'h0/* 0*/ : T339;
    dramBank4PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T349;
    dramBank4_ready_received <= reset ? 1'h0/* 0*/ : T353;
    dramBank3_valid_received_7 <= reset ? 1'h0/* 0*/ : T369;
    dramBank3_valid_received_6 <= reset ? 1'h0/* 0*/ : T380;
    dramBank3_valid_received_5 <= reset ? 1'h0/* 0*/ : T390;
    dramBank3_valid_received_4 <= reset ? 1'h0/* 0*/ : T400;
    dramBank3_valid_received_3 <= reset ? 1'h0/* 0*/ : T410;
    dramBank3_valid_received_2 <= reset ? 1'h0/* 0*/ : T420;
    dramBank3_valid_received_1 <= reset ? 1'h0/* 0*/ : T430;
    dramBank3_valid_received_0 <= reset ? 1'h0/* 0*/ : T439;
    dramBank3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T449;
    dramBank3_ready_received <= reset ? 1'h0/* 0*/ : T453;
    dramBank2_valid_received_7 <= reset ? 1'h0/* 0*/ : T469;
    dramBank2_valid_received_6 <= reset ? 1'h0/* 0*/ : T480;
    dramBank2_valid_received_5 <= reset ? 1'h0/* 0*/ : T490;
    dramBank2_valid_received_4 <= reset ? 1'h0/* 0*/ : T500;
    dramBank2_valid_received_3 <= reset ? 1'h0/* 0*/ : T510;
    dramBank2_valid_received_2 <= reset ? 1'h0/* 0*/ : T520;
    dramBank2_valid_received_1 <= reset ? 1'h0/* 0*/ : T530;
    dramBank2_valid_received_0 <= reset ? 1'h0/* 0*/ : T539;
    dramBank2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T549;
    dramBank2_ready_received <= reset ? 1'h0/* 0*/ : T553;
    dramBank1_valid_received_7 <= reset ? 1'h0/* 0*/ : T569;
    dramBank1_valid_received_6 <= reset ? 1'h0/* 0*/ : T580;
    dramBank1_valid_received_5 <= reset ? 1'h0/* 0*/ : T590;
    dramBank1_valid_received_4 <= reset ? 1'h0/* 0*/ : T600;
    dramBank1_valid_received_3 <= reset ? 1'h0/* 0*/ : T610;
    dramBank1_valid_received_2 <= reset ? 1'h0/* 0*/ : T620;
    dramBank1_valid_received_1 <= reset ? 1'h0/* 0*/ : T630;
    dramBank1_valid_received_0 <= reset ? 1'h0/* 0*/ : T639;
    dramBank1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T649;
    dramBank1_ready_received <= reset ? 1'h0/* 0*/ : T653;
    dramBank0_valid_received_7 <= reset ? 1'h0/* 0*/ : T668;
    dramBank0_valid_received_6 <= reset ? 1'h0/* 0*/ : T679;
    dramBank0_valid_received_5 <= reset ? 1'h0/* 0*/ : T689;
    dramBank0_valid_received_4 <= reset ? 1'h0/* 0*/ : T699;
    dramBank0_valid_received_3 <= reset ? 1'h0/* 0*/ : T709;
    dramBank0_valid_received_2 <= reset ? 1'h0/* 0*/ : T719;
    dramBank0_valid_received_1 <= reset ? 1'h0/* 0*/ : T729;
    dramBank0_valid_received_0 <= reset ? 1'h0/* 0*/ : T738;
    dramBank0PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T748;
    dramBank0_ready_received <= reset ? 1'h0/* 0*/ : T752;
    subStateTh_6 <= reset ? 1'h0/* 0*/ : T756;
    if(reset) begin
      State_6 <= 8'h0/* 0*/;
    end else if(T762) begin
      State_6 <= T2240;
    end
    if(reset) begin
      State_5 <= 8'h0/* 0*/;
    end else if(T778) begin
      State_5 <= T1508;
    end
    if(T839) begin
      inputReg_7_addr <= T845;
    end
    if(T849) begin
      inputReg_6_addr <= T851;
    end
    if(T855) begin
      inputReg_5_addr <= T857;
    end
    if(T862) begin
      inputReg_4_addr <= T864;
    end
    if(T869) begin
      inputReg_3_addr <= T871;
    end
    if(T876) begin
      inputReg_2_addr <= T878;
    end
    if(T883) begin
      inputReg_1_addr <= T885;
    end
    if(T889) begin
      inputReg_0_addr <= T891;
    end
    if(reset) begin
      rb7RowAddr_7 <= 32'h0/* 0*/;
    end else if(T935) begin
      rb7RowAddr_7 <= T937;
    end
    if(reset) begin
      rb7RowAddr_6 <= 32'h0/* 0*/;
    end else if(T943) begin
      rb7RowAddr_6 <= T945;
    end
    if(reset) begin
      rb7RowAddr_5 <= 32'h0/* 0*/;
    end else if(T951) begin
      rb7RowAddr_5 <= T952;
    end
    if(reset) begin
      rb7RowAddr_4 <= 32'h0/* 0*/;
    end else if(T958) begin
      rb7RowAddr_4 <= T960;
    end
    if(reset) begin
      rb7RowAddr_3 <= 32'h0/* 0*/;
    end else if(T966) begin
      rb7RowAddr_3 <= T968;
    end
    if(reset) begin
      rb7RowAddr_2 <= 32'h0/* 0*/;
    end else if(T974) begin
      rb7RowAddr_2 <= T976;
    end
    if(reset) begin
      rb7RowAddr_1 <= 32'h0/* 0*/;
    end else if(T982) begin
      rb7RowAddr_1 <= T984;
    end
    if(reset) begin
      rb7RowAddr_0 <= 32'h0/* 0*/;
    end else if(T989) begin
      rb7RowAddr_0 <= T991;
    end
    if(reset) begin
      rb6RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1007) begin
      rb6RowAddr_7 <= T1009;
    end
    if(reset) begin
      rb6RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1015) begin
      rb6RowAddr_6 <= T1017;
    end
    if(reset) begin
      rb6RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1023) begin
      rb6RowAddr_5 <= T1024;
    end
    if(reset) begin
      rb6RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1030) begin
      rb6RowAddr_4 <= T1032;
    end
    if(reset) begin
      rb6RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1038) begin
      rb6RowAddr_3 <= T1040;
    end
    if(reset) begin
      rb6RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1046) begin
      rb6RowAddr_2 <= T1048;
    end
    if(reset) begin
      rb6RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1054) begin
      rb6RowAddr_1 <= T1056;
    end
    if(reset) begin
      rb6RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1061) begin
      rb6RowAddr_0 <= T1063;
    end
    if(reset) begin
      rb5RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1079) begin
      rb5RowAddr_7 <= T1081;
    end
    if(reset) begin
      rb5RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1087) begin
      rb5RowAddr_6 <= T1089;
    end
    if(reset) begin
      rb5RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1095) begin
      rb5RowAddr_5 <= T1096;
    end
    if(reset) begin
      rb5RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1102) begin
      rb5RowAddr_4 <= T1104;
    end
    if(reset) begin
      rb5RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1110) begin
      rb5RowAddr_3 <= T1112;
    end
    if(reset) begin
      rb5RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1118) begin
      rb5RowAddr_2 <= T1120;
    end
    if(reset) begin
      rb5RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1126) begin
      rb5RowAddr_1 <= T1128;
    end
    if(reset) begin
      rb5RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1133) begin
      rb5RowAddr_0 <= T1135;
    end
    if(reset) begin
      rb4RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1151) begin
      rb4RowAddr_7 <= T1153;
    end
    if(reset) begin
      rb4RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1159) begin
      rb4RowAddr_6 <= T1161;
    end
    if(reset) begin
      rb4RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1167) begin
      rb4RowAddr_5 <= T1168;
    end
    if(reset) begin
      rb4RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1174) begin
      rb4RowAddr_4 <= T1176;
    end
    if(reset) begin
      rb4RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1182) begin
      rb4RowAddr_3 <= T1184;
    end
    if(reset) begin
      rb4RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1190) begin
      rb4RowAddr_2 <= T1192;
    end
    if(reset) begin
      rb4RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1198) begin
      rb4RowAddr_1 <= T1200;
    end
    if(reset) begin
      rb4RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1205) begin
      rb4RowAddr_0 <= T1207;
    end
    if(reset) begin
      rb3RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1223) begin
      rb3RowAddr_7 <= T1225;
    end
    if(reset) begin
      rb3RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1231) begin
      rb3RowAddr_6 <= T1233;
    end
    if(reset) begin
      rb3RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1239) begin
      rb3RowAddr_5 <= T1240;
    end
    if(reset) begin
      rb3RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1246) begin
      rb3RowAddr_4 <= T1248;
    end
    if(reset) begin
      rb3RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1254) begin
      rb3RowAddr_3 <= T1256;
    end
    if(reset) begin
      rb3RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1262) begin
      rb3RowAddr_2 <= T1264;
    end
    if(reset) begin
      rb3RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1270) begin
      rb3RowAddr_1 <= T1272;
    end
    if(reset) begin
      rb3RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1277) begin
      rb3RowAddr_0 <= T1279;
    end
    if(reset) begin
      rb2RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1295) begin
      rb2RowAddr_7 <= T1297;
    end
    if(reset) begin
      rb2RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1303) begin
      rb2RowAddr_6 <= T1305;
    end
    if(reset) begin
      rb2RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1311) begin
      rb2RowAddr_5 <= T1312;
    end
    if(reset) begin
      rb2RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1318) begin
      rb2RowAddr_4 <= T1320;
    end
    if(reset) begin
      rb2RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1326) begin
      rb2RowAddr_3 <= T1328;
    end
    if(reset) begin
      rb2RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1334) begin
      rb2RowAddr_2 <= T1336;
    end
    if(reset) begin
      rb2RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1342) begin
      rb2RowAddr_1 <= T1344;
    end
    if(reset) begin
      rb2RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1349) begin
      rb2RowAddr_0 <= T1351;
    end
    if(reset) begin
      rb1RowAddr_7 <= 32'h0/* 0*/;
    end else if(T1367) begin
      rb1RowAddr_7 <= T1369;
    end
    if(reset) begin
      rb1RowAddr_6 <= 32'h0/* 0*/;
    end else if(T1375) begin
      rb1RowAddr_6 <= T1377;
    end
    if(reset) begin
      rb1RowAddr_5 <= 32'h0/* 0*/;
    end else if(T1383) begin
      rb1RowAddr_5 <= T1384;
    end
    if(reset) begin
      rb1RowAddr_4 <= 32'h0/* 0*/;
    end else if(T1390) begin
      rb1RowAddr_4 <= T1392;
    end
    if(reset) begin
      rb1RowAddr_3 <= 32'h0/* 0*/;
    end else if(T1398) begin
      rb1RowAddr_3 <= T1400;
    end
    if(reset) begin
      rb1RowAddr_2 <= 32'h0/* 0*/;
    end else if(T1406) begin
      rb1RowAddr_2 <= T1408;
    end
    if(reset) begin
      rb1RowAddr_1 <= 32'h0/* 0*/;
    end else if(T1414) begin
      rb1RowAddr_1 <= T1416;
    end
    if(reset) begin
      rb1RowAddr_0 <= 32'h0/* 0*/;
    end else if(T1421) begin
      rb1RowAddr_0 <= T1423;
    end
    if(reset) begin
      rb0RowAddr_7 <= 32'h1/* 1*/;
    end else if(T1439) begin
      rb0RowAddr_7 <= T1441;
    end
    if(reset) begin
      rb0RowAddr_6 <= 32'h1/* 1*/;
    end else if(T1447) begin
      rb0RowAddr_6 <= T1449;
    end
    if(reset) begin
      rb0RowAddr_5 <= 32'h1/* 1*/;
    end else if(T1455) begin
      rb0RowAddr_5 <= T1456;
    end
    if(reset) begin
      rb0RowAddr_4 <= 32'h1/* 1*/;
    end else if(T1462) begin
      rb0RowAddr_4 <= T1464;
    end
    if(reset) begin
      rb0RowAddr_3 <= 32'h1/* 1*/;
    end else if(T1470) begin
      rb0RowAddr_3 <= T1472;
    end
    if(reset) begin
      rb0RowAddr_2 <= 32'h1/* 1*/;
    end else if(T1478) begin
      rb0RowAddr_2 <= T1480;
    end
    if(reset) begin
      rb0RowAddr_1 <= 32'h1/* 1*/;
    end else if(T1486) begin
      rb0RowAddr_1 <= T1488;
    end
    if(reset) begin
      rb0RowAddr_0 <= 32'h1/* 1*/;
    end else if(T1493) begin
      rb0RowAddr_0 <= T1495;
    end
    if(reset) begin
      EmitReturnState_7 <= 8'h0/* 0*/;
    end else if(T1532) begin
      EmitReturnState_7 <= T1548;
    end
    if(reset) begin
      EmitReturnState_6 <= 8'h0/* 0*/;
    end else if(T1560) begin
      EmitReturnState_6 <= T1576;
    end
    if(reset) begin
      EmitReturnState_5 <= 8'h0/* 0*/;
    end else if(T1588) begin
      EmitReturnState_5 <= T1596;
    end
    if(reset) begin
      EmitReturnState_4 <= 8'h0/* 0*/;
    end else if(T1608) begin
      EmitReturnState_4 <= T1625;
    end
    if(reset) begin
      EmitReturnState_3 <= 8'h0/* 0*/;
    end else if(T1637) begin
      EmitReturnState_3 <= T1654;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T1666) begin
      EmitReturnState_2 <= T1683;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T1695) begin
      EmitReturnState_1 <= T1712;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T1723) begin
      EmitReturnState_0 <= T1740;
    end
    if(reset) begin
      State_4 <= 8'h0/* 0*/;
    end else if(T1777) begin
      State_4 <= T1814;
    end
    if(reset) begin
      State_3 <= 8'h0/* 0*/;
    end else if(T1863) begin
      State_3 <= T1900;
    end
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T1949) begin
      State_2 <= T1986;
    end
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T2035) begin
      State_1 <= T2072;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T2120) begin
      State_0 <= T2157;
    end
    subStateTh_5 <= reset ? 1'h0/* 0*/ : T2292;
    subStateTh_4 <= reset ? 1'h0/* 0*/ : T2304;
    subStateTh_3 <= reset ? 1'h0/* 0*/ : T2316;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T2328;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T2340;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T2352;
    dramBank7_valid_received_7 <= reset ? 1'h0/* 0*/ : T2389;
    dramBank7_valid_received_6 <= reset ? 1'h0/* 0*/ : T2400;
    dramBank7_valid_received_5 <= reset ? 1'h0/* 0*/ : T2410;
    dramBank7_valid_received_4 <= reset ? 1'h0/* 0*/ : T2420;
    dramBank7_valid_received_3 <= reset ? 1'h0/* 0*/ : T2430;
    dramBank7_valid_received_2 <= reset ? 1'h0/* 0*/ : T2440;
    dramBank7_valid_received_1 <= reset ? 1'h0/* 0*/ : T2450;
    dramBank7_valid_received_0 <= reset ? 1'h0/* 0*/ : T2459;
    dramBank6PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2480;
    dramBank5PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2495;
    dramBank4PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2510;
    dramBank3PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2525;
    dramBank2PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2540;
    dramBank1PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2555;
    dramBank0PortHadValidRequest_7 <= reset ? 1'h0/* 0*/ : T2569;
    dramBank7PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2586;
    dramBank6PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2601;
    dramBank5PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2616;
    dramBank4PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2631;
    dramBank3PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2646;
    dramBank2PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2661;
    dramBank1PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2676;
    dramBank0PortHadValidRequest_6 <= reset ? 1'h0/* 0*/ : T2690;
    dramBank7PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2707;
    dramBank6PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2722;
    dramBank5PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2737;
    dramBank4PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2752;
    dramBank3PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2767;
    dramBank2PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2782;
    dramBank1PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2797;
    dramBank0PortHadValidRequest_5 <= reset ? 1'h0/* 0*/ : T2811;
    dramBank7PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2828;
    dramBank6PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2843;
    dramBank5PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2858;
    dramBank4PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2873;
    dramBank3PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2888;
    dramBank2PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2903;
    dramBank1PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2918;
    dramBank0PortHadValidRequest_4 <= reset ? 1'h0/* 0*/ : T2932;
    dramBank7PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2949;
    dramBank6PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2964;
    dramBank5PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2979;
    dramBank4PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T2994;
    dramBank3PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3009;
    dramBank2PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3024;
    dramBank1PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3039;
    dramBank0PortHadValidRequest_3 <= reset ? 1'h0/* 0*/ : T3053;
    dramBank7PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3070;
    dramBank6PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3085;
    dramBank5PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3100;
    dramBank4PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3115;
    dramBank3PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3130;
    dramBank2PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3145;
    dramBank1PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3160;
    dramBank0PortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T3174;
    dramBank7PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3191;
    dramBank6PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3206;
    dramBank5PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3221;
    dramBank4PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3236;
    dramBank3PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3251;
    dramBank2PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3266;
    dramBank1PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3281;
    dramBank0PortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T3295;
    dramBank7PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3312;
    dramBank6PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3327;
    dramBank5PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3342;
    dramBank4PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3357;
    dramBank3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3372;
    dramBank2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3387;
    dramBank1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3402;
    dramBank0PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T3416;
    if(T839) begin
      inputTag_7 <= T3538;
    end
    if(T849) begin
      inputTag_6 <= T3542;
    end
    if(T855) begin
      inputTag_5 <= T3546;
    end
    if(T862) begin
      inputTag_4 <= T3550;
    end
    if(T869) begin
      inputTag_3 <= T3554;
    end
    if(T876) begin
      inputTag_2 <= T3558;
    end
    if(T883) begin
      inputTag_1 <= T3562;
    end
    if(T889) begin
      inputTag_0 <= T3565;
    end
  end
endmodule

module RREncode_62(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_63(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_64(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_62 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_63 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_64 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_23(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank1_req_ready,
    output mainOff_dramBank1_req_valid,
    output[31:0] mainOff_dramBank1_req_bits,
    output[9:0] mainOff_dramBank1_req_tag,
    output mainOff_dramBank1_rep_ready,
    input  mainOff_dramBank1_rep_valid,
    input [31:0] mainOff_dramBank1_rep_bits,
    input [9:0] mainOff_dramBank1_rep_tag,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire mainComp_mainOff_dramBank1_rep_ready;
  wire mainComp_mainOff_dramBank1_req_valid;
  wire[9:0] mainComp_mainOff_dramBank1_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank0_rep_ready;
  wire mainComp_mainOff_dramBank0_req_valid;
  wire[9:0] mainComp_mainOff_dramBank0_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank2_rep_ready = mainComp_mainOff_dramBank2_rep_ready;
  assign mainOff_dramBank2_req_valid = mainComp_mainOff_dramBank2_req_valid;
  assign mainOff_dramBank2_req_tag = mainComp_mainOff_dramBank2_req_tag;
  assign mainOff_dramBank1_rep_ready = mainComp_mainOff_dramBank1_rep_ready;
  assign mainOff_dramBank1_req_valid = mainComp_mainOff_dramBank1_req_valid;
  assign mainOff_dramBank1_req_tag = mainComp_mainOff_dramBank1_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  dram_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank0_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank0_req_valid( mainComp_mainOff_dramBank0_req_valid ),
       .mainOff_dramBank0_req_bits(  ),
       .mainOff_dramBank0_req_tag( mainComp_mainOff_dramBank0_req_tag ),
       .mainOff_dramBank0_rep_ready( mainComp_mainOff_dramBank0_rep_ready ),
       .mainOff_dramBank0_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank0_rep_bits(  ),
       .mainOff_dramBank0_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank1_req_ready( mainOff_dramBank1_req_ready ),
       .mainOff_dramBank1_req_valid( mainComp_mainOff_dramBank1_req_valid ),
       .mainOff_dramBank1_req_bits(  ),
       .mainOff_dramBank1_req_tag( mainComp_mainOff_dramBank1_req_tag ),
       .mainOff_dramBank1_rep_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .mainOff_dramBank1_rep_valid( mainOff_dramBank1_rep_valid ),
       .mainOff_dramBank1_rep_bits(  ),
       .mainOff_dramBank1_rep_tag( mainOff_dramBank1_rep_tag ),
       .mainOff_dramBank2_req_ready( mainOff_dramBank2_req_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( mainOff_dramBank2_rep_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( mainOff_dramBank2_rep_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_8 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank0_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank0_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank0_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_65(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_66(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_67(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_65 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_66 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_67 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_24(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank2_req_ready,
    output mainOff_dramBank2_req_valid,
    output[31:0] mainOff_dramBank2_req_bits,
    output[9:0] mainOff_dramBank2_req_tag,
    output mainOff_dramBank2_rep_ready,
    input  mainOff_dramBank2_rep_valid,
    input [31:0] mainOff_dramBank2_rep_bits,
    input [9:0] mainOff_dramBank2_rep_tag,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank1_rep_ready;
  wire mainComp_mainOff_dramBank1_req_valid;
  wire[9:0] mainComp_mainOff_dramBank1_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank2_rep_ready = mainComp_mainOff_dramBank2_rep_ready;
  assign mainOff_dramBank2_req_valid = mainComp_mainOff_dramBank2_req_valid;
  assign mainOff_dramBank2_req_tag = mainComp_mainOff_dramBank2_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_23 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank1_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank1_req_valid( mainComp_mainOff_dramBank1_req_valid ),
       .mainOff_dramBank1_req_bits(  ),
       .mainOff_dramBank1_req_tag( mainComp_mainOff_dramBank1_req_tag ),
       .mainOff_dramBank1_rep_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .mainOff_dramBank1_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank1_rep_bits(  ),
       .mainOff_dramBank1_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank2_req_ready( mainOff_dramBank2_req_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( mainOff_dramBank2_rep_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( mainOff_dramBank2_rep_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_9 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank1_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank1_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_68(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_69(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_70(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_68 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_69 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_70 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_25(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank3_req_ready,
    output mainOff_dramBank3_req_valid,
    output[31:0] mainOff_dramBank3_req_bits,
    output[9:0] mainOff_dramBank3_req_tag,
    output mainOff_dramBank3_rep_ready,
    input  mainOff_dramBank3_rep_valid,
    input [31:0] mainOff_dramBank3_rep_bits,
    input [9:0] mainOff_dramBank3_rep_tag,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank2_rep_ready;
  wire mainComp_mainOff_dramBank2_req_valid;
  wire[9:0] mainComp_mainOff_dramBank2_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank3_rep_ready = mainComp_mainOff_dramBank3_rep_ready;
  assign mainOff_dramBank3_req_valid = mainComp_mainOff_dramBank3_req_valid;
  assign mainOff_dramBank3_req_tag = mainComp_mainOff_dramBank3_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_24 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank2_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank2_req_valid( mainComp_mainOff_dramBank2_req_valid ),
       .mainOff_dramBank2_req_bits(  ),
       .mainOff_dramBank2_req_tag( mainComp_mainOff_dramBank2_req_tag ),
       .mainOff_dramBank2_rep_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .mainOff_dramBank2_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank2_rep_bits(  ),
       .mainOff_dramBank2_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank3_req_ready( mainOff_dramBank3_req_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( mainOff_dramBank3_rep_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( mainOff_dramBank3_rep_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_10 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank2_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank2_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_71(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_72(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_73(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_71 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_72 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_73 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_26(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank4_req_ready,
    output mainOff_dramBank4_req_valid,
    output[31:0] mainOff_dramBank4_req_bits,
    output[9:0] mainOff_dramBank4_req_tag,
    output mainOff_dramBank4_rep_ready,
    input  mainOff_dramBank4_rep_valid,
    input [31:0] mainOff_dramBank4_rep_bits,
    input [9:0] mainOff_dramBank4_rep_tag,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank3_rep_ready;
  wire mainComp_mainOff_dramBank3_req_valid;
  wire[9:0] mainComp_mainOff_dramBank3_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank4_rep_ready = mainComp_mainOff_dramBank4_rep_ready;
  assign mainOff_dramBank4_req_valid = mainComp_mainOff_dramBank4_req_valid;
  assign mainOff_dramBank4_req_tag = mainComp_mainOff_dramBank4_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_25 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank3_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank3_req_valid( mainComp_mainOff_dramBank3_req_valid ),
       .mainOff_dramBank3_req_bits(  ),
       .mainOff_dramBank3_req_tag( mainComp_mainOff_dramBank3_req_tag ),
       .mainOff_dramBank3_rep_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .mainOff_dramBank3_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank3_rep_bits(  ),
       .mainOff_dramBank3_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank4_req_ready( mainOff_dramBank4_req_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( mainOff_dramBank4_rep_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( mainOff_dramBank4_rep_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_11 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank3_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank3_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_74(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_75(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_76(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_74 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_75 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_76 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_27(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank5_req_ready,
    output mainOff_dramBank5_req_valid,
    output[31:0] mainOff_dramBank5_req_bits,
    output[9:0] mainOff_dramBank5_req_tag,
    output mainOff_dramBank5_rep_ready,
    input  mainOff_dramBank5_rep_valid,
    input [31:0] mainOff_dramBank5_rep_bits,
    input [9:0] mainOff_dramBank5_rep_tag,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank4_rep_ready;
  wire mainComp_mainOff_dramBank4_req_valid;
  wire[9:0] mainComp_mainOff_dramBank4_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank5_rep_ready = mainComp_mainOff_dramBank5_rep_ready;
  assign mainOff_dramBank5_req_valid = mainComp_mainOff_dramBank5_req_valid;
  assign mainOff_dramBank5_req_tag = mainComp_mainOff_dramBank5_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_26 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank4_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank4_req_valid( mainComp_mainOff_dramBank4_req_valid ),
       .mainOff_dramBank4_req_bits(  ),
       .mainOff_dramBank4_req_tag( mainComp_mainOff_dramBank4_req_tag ),
       .mainOff_dramBank4_rep_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .mainOff_dramBank4_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank4_rep_bits(  ),
       .mainOff_dramBank4_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank5_req_ready( mainOff_dramBank5_req_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( mainOff_dramBank5_rep_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( mainOff_dramBank5_rep_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_12 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank4_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank4_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank4_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_77(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_78(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_79(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_77 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_78 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_79 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_28(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank6_req_ready,
    output mainOff_dramBank6_req_valid,
    output[31:0] mainOff_dramBank6_req_bits,
    output[9:0] mainOff_dramBank6_req_tag,
    output mainOff_dramBank6_rep_ready,
    input  mainOff_dramBank6_rep_valid,
    input [31:0] mainOff_dramBank6_rep_bits,
    input [9:0] mainOff_dramBank6_rep_tag,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank5_rep_ready;
  wire mainComp_mainOff_dramBank5_req_valid;
  wire[9:0] mainComp_mainOff_dramBank5_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank6_rep_ready = mainComp_mainOff_dramBank6_rep_ready;
  assign mainOff_dramBank6_req_valid = mainComp_mainOff_dramBank6_req_valid;
  assign mainOff_dramBank6_req_tag = mainComp_mainOff_dramBank6_req_tag;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_27 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank5_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank5_req_valid( mainComp_mainOff_dramBank5_req_valid ),
       .mainOff_dramBank5_req_bits(  ),
       .mainOff_dramBank5_req_tag( mainComp_mainOff_dramBank5_req_tag ),
       .mainOff_dramBank5_rep_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .mainOff_dramBank5_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank5_rep_bits(  ),
       .mainOff_dramBank5_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank6_req_ready( mainOff_dramBank6_req_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( mainOff_dramBank6_rep_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( mainOff_dramBank6_rep_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_13 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank5_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank5_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank5_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_80(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_81(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_82(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[7:0] State_0;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[31:0] T28;
  wire[31:0] T29;
  reg[31:0] counter_0;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[7:0] T39;
  wire T40;
  wire[31:0] T41;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire sThreadEncoder_io_chosen;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire AllOffloadsReady;
  reg[9:0] inputTag_0;
  wire[9:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T11 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T10 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T10 = subStateTh_0 == 1'h1/* 1*/;
  assign T11 = T73 && T12;
  assign T12 = State_0 != 8'hff/* 255*/;
  assign T13 = T24 || T14;
  assign T14 = T18 && T15;
  assign T15 = T16;
  assign T16 = T17[1'h0/* 0*/:1'h0/* 0*/];
  assign T17 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T18 = T23 && T19;
  assign T19 = T21 == T20;
  assign T20 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T21 = State_0 & T22;
  assign T22 = {4'h8/* 8*/{T15}};
  assign T23 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T24 = T44 || T25;
  assign T25 = T26 && T15;
  assign T26 = T32 && T27;
  assign T27 = T28 == 32'h0/* 0*/;
  assign T28 = counter_0 & T29;
  assign T29 = {6'h20/* 32*/{T15}};
  assign T30 = T36 || T31;
  assign T31 = T32 && T15;
  assign T32 = T35 && T33;
  assign T33 = T21 == T34;
  assign T34 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T35 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T36 = T37 && T15;
  assign T37 = T40 && T38;
  assign T38 = T21 == T39;
  assign T39 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T41 = T31 ? T43 : T42;
  assign T42 = T36 ? 32'ha/* 10*/ : counter_0;
  assign T43 = T28 - 32'h1/* 1*/;
  assign T44 = T45 || T36;
  assign T45 = T53 || T46;
  assign T46 = T47 && T2;
  assign T47 = T48 && io_out_ready;
  assign T48 = T52 && T49;
  assign T49 = T50 == 8'hff/* 255*/;
  assign T50 = State_0 & T51;
  assign T51 = {4'h8/* 8*/{T2}};
  assign T52 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T53 = T60 && T54;
  assign T54 = T55;
  assign T55 = T56[1'h0/* 0*/:1'h0/* 0*/];
  assign T56 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T57 = T59 && T58;
  assign T58 = State_0 == 8'h0/* 0*/;
  assign T59 = subStateTh_0 == 1'h0/* 0*/;
  assign T60 = T61 && io_in_valid;
  assign T61 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T62 = T14 ? 8'hff/* 255*/ : T63;
  assign T63 = T25 ? T72 : T64;
  assign T64 = T36 ? T71 : T65;
  assign T65 = T46 ? T68 : T66;
  assign T66 = T53 ? T67 : State_0;
  assign T67 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T68 = EmitReturnState_0 & T69;
  assign T69 = {4'h8/* 8*/{T2}};
  assign T70 = T14 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T71 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T72 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T73 = T75 && T74;
  assign T74 = State_0 != 8'h0/* 0*/;
  assign T75 = AllOffloadsReady && T76;
  assign T76 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T77 = T53 ? io_in_tag : inputTag_0;
  assign io_out_valid = T78;
  assign T78 = T80 && T79;
  assign T79 = T50 == 8'hff/* 255*/;
  assign T80 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T81;
  assign T81 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_80 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_81 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_82 sThreadEncoder(
       .io_valid_0( T57 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T13) begin
      State_0 <= T62;
    end
    if(T30) begin
      counter_0 <= T41;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T14) begin
      EmitReturnState_0 <= T70;
    end
    if(T53) begin
      inputTag_0 <= T77;
    end
  end
endmodule

module gOffloadedComponent_29(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_dramBank7_req_ready,
    output mainOff_dramBank7_req_valid,
    output[31:0] mainOff_dramBank7_req_bits,
    output[9:0] mainOff_dramBank7_req_tag,
    output mainOff_dramBank7_rep_ready,
    input  mainOff_dramBank7_rep_valid,
    input [31:0] mainOff_dramBank7_rep_bits,
    input [9:0] mainOff_dramBank7_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_dramBank6_rep_ready;
  wire mainComp_mainOff_dramBank6_req_valid;
  wire[9:0] mainComp_mainOff_dramBank6_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_dramBank7_rep_ready = mainComp_mainOff_dramBank7_rep_ready;
  assign mainOff_dramBank7_req_valid = mainComp_mainOff_dramBank7_req_valid;
  assign mainOff_dramBank7_req_tag = mainComp_mainOff_dramBank7_req_tag;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_28 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank6_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank6_req_valid( mainComp_mainOff_dramBank6_req_valid ),
       .mainOff_dramBank6_req_bits(  ),
       .mainOff_dramBank6_req_tag( mainComp_mainOff_dramBank6_req_tag ),
       .mainOff_dramBank6_rep_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .mainOff_dramBank6_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank6_rep_bits(  ),
       .mainOff_dramBank6_rep_tag( offComp_io_out_tag ),
       .mainOff_dramBank7_req_ready( mainOff_dramBank7_req_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( mainOff_dramBank7_rep_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( mainOff_dramBank7_rep_tag ));
  dramBank_14 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank6_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank6_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank6_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_83(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_84(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_85(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module dramBank_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire T0;
  wire sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_0;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  wire vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_0;
  wire T9;
  reg[0:0] subStateTh_0;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire rThreadEncoder_io_chosen;
  wire T19;
  wire AllOffloadsReady;
  wire T20;
  wire T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire[31:0] T31;
  reg[31:0] counter_0;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[7:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[7:0] T41;
  wire T42;
  wire[31:0] T43;
  wire[31:0] T44;
  wire[31:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire T75;
  wire[9:0] T76;
  wire[9:0] T77;
  reg[9:0] inputTag_0;
  wire[9:0] T78;
  wire T79;
  wire T80;
  wire T81;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T1 = T75 && T2;
  assign T2 = State_0 == 8'h0/* 0*/;
  assign T3 = T26 || T4;
  assign T4 = T20 && T5;
  assign T5 = T6;
  assign T6 = T7[1'h0/* 0*/:1'h0/* 0*/];
  assign T7 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T9 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T9 = subStateTh_0 == 1'h1/* 1*/;
  assign T10 = T13 ? 1'h1/* 1*/ : T11;
  assign T11 = T12 ? 1'h0/* 0*/ : subStateTh_0;
  assign T12 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T13 = T15 && T14;
  assign T14 = State_0 != 8'hff/* 255*/;
  assign T15 = T17 && T16;
  assign T16 = State_0 != 8'h0/* 0*/;
  assign T17 = AllOffloadsReady && T18;
  assign T18 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign T19 = subStateTh_0 == 1'h0/* 0*/;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T20 = T25 && T21;
  assign T21 = T23 == T22;
  assign T22 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T23 = State_0 & T24;
  assign T24 = {4'h8/* 8*/{T5}};
  assign T25 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T26 = T46 || T27;
  assign T27 = T28 && T5;
  assign T28 = T34 && T29;
  assign T29 = T30 == 32'h0/* 0*/;
  assign T30 = counter_0 & T31;
  assign T31 = {6'h20/* 32*/{T5}};
  assign T32 = T38 || T33;
  assign T33 = T34 && T5;
  assign T34 = T37 && T35;
  assign T35 = T23 == T36;
  assign T36 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T37 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T38 = T39 && T5;
  assign T39 = T42 && T40;
  assign T40 = T23 == T41;
  assign T41 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T42 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T43 = T33 ? T45 : T44;
  assign T44 = T38 ? 32'ha/* 10*/ : counter_0;
  assign T45 = T30 - 32'h1/* 1*/;
  assign T46 = T47 || T38;
  assign T47 = T58 || T48;
  assign T48 = T52 && T49;
  assign T49 = T50;
  assign T50 = T51[1'h0/* 0*/:1'h0/* 0*/];
  assign T51 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T52 = T53 && io_out_ready;
  assign T53 = T57 && T54;
  assign T54 = T55 == 8'hff/* 255*/;
  assign T55 = State_0 & T56;
  assign T56 = {4'h8/* 8*/{T49}};
  assign T57 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T58 = T62 && T59;
  assign T59 = T60;
  assign T60 = T61[1'h0/* 0*/:1'h0/* 0*/];
  assign T61 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T62 = T63 && io_in_valid;
  assign T63 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T64 = T4 ? 8'hff/* 255*/ : T65;
  assign T65 = T27 ? T74 : T66;
  assign T66 = T38 ? T73 : T67;
  assign T67 = T48 ? T70 : T68;
  assign T68 = T58 ? T69 : State_0;
  assign T69 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T70 = EmitReturnState_0 & T71;
  assign T71 = {4'h8/* 8*/{T49}};
  assign T72 = T4 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T73 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T74 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign io_out_tag = T76;
  assign T76 = inputTag_0 & T77;
  assign T77 = {4'ha/* 10*/{T49}};
  assign T78 = T58 ? io_in_tag : inputTag_0;
  assign io_out_valid = T79;
  assign T79 = T81 && T80;
  assign T80 = T55 == 8'hff/* 255*/;
  assign T81 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_83 rThreadEncoder(
       .io_valid_0( T19 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_84 vThreadEncoder(
       .io_valid_0( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_85 sThreadEncoder(
       .io_valid_0( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_0 <= T64;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T10;
    if(T32) begin
      counter_0 <= T43;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_0 <= T72;
    end
    if(T58) begin
      inputTag_0 <= T78;
    end
  end
endmodule

module gOffloadedComponent_30(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_dramBank7_rep_ready;
  wire mainComp_mainOff_dramBank7_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_dramBank7_req_tag;
  wire offComp_io_out_valid;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_29 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dramBank7_req_ready( offComp_io_in_ready ),
       .mainOff_dramBank7_req_valid( mainComp_mainOff_dramBank7_req_valid ),
       .mainOff_dramBank7_req_bits(  ),
       .mainOff_dramBank7_req_tag( mainComp_mainOff_dramBank7_req_tag ),
       .mainOff_dramBank7_rep_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .mainOff_dramBank7_rep_valid( offComp_io_out_valid ),
       .mainOff_dramBank7_rep_bits(  ),
       .mainOff_dramBank7_rep_tag( offComp_io_out_tag ));
  dramBank_15 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dramBank7_req_valid ),
       .io_in_bits(  ),
       .io_in_tag( mainComp_mainOff_dramBank7_req_tag ),
       .io_out_ready( mainComp_mainOff_dramBank7_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_31(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_dram_req_valid;
  wire[31:0] mainComp_mainOff_dram_req_bits_addr;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[127:0] mainComp_io_out_bits_data;
  wire mainComp_mainOff_dram_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_dram_req_tag;
  wire offComp_io_out_valid;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_bits_data = mainComp_io_out_bits_data;
  gOffloadedComponent_22 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_data( mainComp_io_out_bits_data ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_dram_req_ready( offComp_io_in_ready ),
       .mainOff_dram_req_valid( mainComp_mainOff_dram_req_valid ),
       .mainOff_dram_req_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .mainOff_dram_req_bits_rw(  ),
       .mainOff_dram_req_bits_cached(  ),
       .mainOff_dram_req_bits_data(  ),
       .mainOff_dram_req_bits_size(  ),
       .mainOff_dram_req_tag( mainComp_mainOff_dram_req_tag ),
       .mainOff_dram_rep_ready( mainComp_mainOff_dram_rep_ready ),
       .mainOff_dram_rep_valid( offComp_io_out_valid ),
       .mainOff_dram_rep_bits_data(  ),
       .mainOff_dram_rep_tag( offComp_io_out_tag ));
  gOffloadedComponent_30 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_dram_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_dram_req_bits_addr ),
       .io_in_bits_rw(  ),
       .io_in_bits_cached(  ),
       .io_in_bits_data(  ),
       .io_in_bits_size(  ),
       .io_in_tag( mainComp_mainOff_dram_req_tag ),
       .io_out_ready( mainComp_mainOff_dram_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_data(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module prMemComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input  io_in_bits_cached,
    input [127:0] io_in_bits_data,
    input [3:0] io_in_bits_size,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[127:0] io_out_bits_data,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] generatedTop_io_out_tag;
  wire generatedTop_io_out_valid;
  wire generatedTop_io_in_ready;
  wire[127:0] generatedTop_io_out_bits_data;

  assign io_out_tag = generatedTop_io_out_tag;
  assign io_out_valid = generatedTop_io_out_valid;
  assign io_in_ready = generatedTop_io_in_ready;
  assign io_out_bits_data = generatedTop_io_out_bits_data;
  gOffloadedComponent_31 generatedTop(.clk(clk), .reset(reset),
       .io_in_ready( generatedTop_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_addr( io_in_bits_addr ),
       .io_in_bits_rw( io_in_bits_rw ),
       .io_in_bits_cached( io_in_bits_cached ),
       .io_in_bits_data( io_in_bits_data ),
       .io_in_bits_size( io_in_bits_size ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( generatedTop_io_out_valid ),
       .io_out_bits_data( generatedTop_io_out_bits_data ),
       .io_out_tag( generatedTop_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_32(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_pageId,
    input [63:0] io_in_bits_rankUpdate,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire[9:0] offComp_io_out_tag;
  wire[3:0] mainComp_mainOff_mem_req_bits_size;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire[127:0] offComp_io_out_bits_data;
  wire[31:0] mainComp_mainOff_mem_req_bits_addr;
  wire mainComp_mainOff_mem_req_valid;
  wire[127:0] mainComp_mainOff_mem_req_bits_data;
  wire mainComp_mainOff_mem_req_bits_cached;
  wire mainComp_mainOff_mem_req_bits_rw;
  wire mainComp_mainOff_mem_rep_ready;
  wire[9:0] mainComp_mainOff_mem_req_tag;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  gOffloadedComponent_21 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_pageId( io_in_bits_pageId ),
       .io_in_bits_rankUpdate( io_in_bits_rankUpdate ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_mem_req_ready( offComp_io_in_ready ),
       .mainOff_mem_req_valid( mainComp_mainOff_mem_req_valid ),
       .mainOff_mem_req_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .mainOff_mem_req_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .mainOff_mem_req_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .mainOff_mem_req_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .mainOff_mem_req_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .mainOff_mem_req_tag( mainComp_mainOff_mem_req_tag ),
       .mainOff_mem_rep_ready( mainComp_mainOff_mem_rep_ready ),
       .mainOff_mem_rep_valid( offComp_io_out_valid ),
       .mainOff_mem_rep_bits_data( offComp_io_out_bits_data ),
       .mainOff_mem_rep_tag( offComp_io_out_tag ));
  prMemComponent_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_mem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_mem_req_bits_rw ),
       .io_in_bits_cached( mainComp_mainOff_mem_req_bits_cached ),
       .io_in_bits_data( mainComp_mainOff_mem_req_bits_data ),
       .io_in_bits_size( mainComp_mainOff_mem_req_bits_size ),
       .io_in_tag( mainComp_mainOff_mem_req_tag ),
       .io_out_ready( mainComp_mainOff_mem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_data( offComp_io_out_bits_data ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gChainedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire source_io_in_ready;
  wire sink_io_in_ready;
  wire source_io_out_valid;
  wire source_io_out_bits_done;
  wire[31:0] source_io_out_bits_pageId;
  wire[9:0] sink_io_out_tag;
  wire[9:0] source_io_out_tag;
  wire sink_io_out_valid;
  wire[63:0] source_io_out_bits_rankUpdate;

  assign io_in_ready = source_io_in_ready;
  assign io_out_tag = sink_io_out_tag;
  assign io_out_valid = sink_io_out_valid;
  gOffloadedComponent_16 source(.clk(clk), .reset(reset),
       .io_in_ready( source_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( sink_io_in_ready ),
       .io_out_valid( source_io_out_valid ),
       .io_out_bits_done( source_io_out_bits_done ),
       .io_out_bits_pageId( source_io_out_bits_pageId ),
       .io_out_bits_rankUpdate( source_io_out_bits_rankUpdate ),
       .io_out_tag( source_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_32 sink(.clk(clk), .reset(reset),
       .io_in_ready( sink_io_in_ready ),
       .io_in_valid( source_io_out_valid ),
       .io_in_bits_done( source_io_out_bits_done ),
       .io_in_bits_pageId( source_io_out_bits_pageId ),
       .io_in_bits_rankUpdate( source_io_out_bits_rankUpdate ),
       .io_in_tag( source_io_out_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( sink_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( sink_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module Top(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_done,
    input [31:0] io_in_bits_startPageId,
    input [31:0] io_in_bits_length,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_done,
    output[31:0] io_out_bits_pageId,
    output[63:0] io_out_bits_rankUpdate,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire generatedTop_io_in_ready;
  wire[9:0] generatedTop_io_out_tag;
  wire generatedTop_io_out_valid;

  assign io_in_ready = generatedTop_io_in_ready;
  assign io_out_tag = generatedTop_io_out_tag;
  assign io_out_valid = generatedTop_io_out_valid;
  gChainedComponent generatedTop(.clk(clk), .reset(reset),
       .io_in_ready( generatedTop_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_done( io_in_bits_done ),
       .io_in_bits_startPageId( io_in_bits_startPageId ),
       .io_in_bits_length( io_in_bits_length ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( generatedTop_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( generatedTop_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

