module RREncode(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_1(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_2(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module KDistribute(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire T0;
  wire sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_0;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  wire vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_0;
  wire T9;
  reg[0:0] subStateTh_0;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire rThreadEncoder_io_chosen;
  wire T19;
  wire AllOffloadsReady;
  wire T20;
  wire T21;
  wire[7:0] T22;
  wire[7:0] T23;
  wire[7:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[7:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire T42;
  wire T43;
  reg[0:0] outputReg_0_pointsFinished;
  wire T44;
  wire T45;
  reg[0:0] inputReg_0_pointsFinished;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  reg[0:0] outputReg_0_centeroidsFinished;
  wire T54;
  wire T55;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  reg[7:0] EmitReturnState_0;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[32:0] T71;
  wire[31:0] T72;
  wire[31:0] T73;
  reg[31:0] broadcastIndex_0;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg[31:0] mode;
  wire T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire[31:0] T86;
  wire[31:0] T87;
  wire[31:0] T88;
  wire[31:0] T89;
  wire[31:0] T90;
  wire[31:0] T91;
  wire[31:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire T102;
  wire[7:0] T103;
  wire T104;
  wire T105;
  wire[9:0] T106;
  wire[9:0] T107;
  reg[9:0] inputTag_0;
  wire[9:0] T108;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T1 = T105 && T2;
  assign T2 = State_0 == 8'h0/* 0*/;
  assign T3 = T26 || T4;
  assign T4 = T20 && T5;
  assign T5 = T6;
  assign T6 = T7[1'h0/* 0*/:1'h0/* 0*/];
  assign T7 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T9 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = 1'h1/* 1*/;
  assign T9 = subStateTh_0 == 1'h1/* 1*/;
  assign T10 = T13 ? 1'h1/* 1*/ : T11;
  assign T11 = T12 ? 1'h0/* 0*/ : subStateTh_0;
  assign T12 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T13 = T15 && T14;
  assign T14 = State_0 != 8'hff/* 255*/;
  assign T15 = T17 && T16;
  assign T16 = State_0 != 8'h0/* 0*/;
  assign T17 = AllOffloadsReady && T18;
  assign T18 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign T19 = subStateTh_0 == 1'h0/* 0*/;
  assign AllOffloadsReady = 1'h1/* 1*/;
  assign T20 = T25 && T21;
  assign T21 = T23 == T22;
  assign T22 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T23 = State_0 & T24;
  assign T24 = {4'h8/* 8*/{T5}};
  assign T25 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T26 = T32 || T27;
  assign T27 = T28 && T5;
  assign T28 = T31 && T29;
  assign T29 = T23 == T30;
  assign T30 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T31 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T32 = T46 || T33;
  assign T33 = T37 && T34;
  assign T34 = T35;
  assign T35 = T36[1'h0/* 0*/:1'h0/* 0*/];
  assign T36 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T37 = T57 && io_out_ready;
  assign io_out_valid = T38;
  assign T38 = T42 && T39;
  assign T39 = T40 == 8'hff/* 255*/;
  assign T40 = State_0 & T41;
  assign T41 = {4'h8/* 8*/{T34}};
  assign T42 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_out_bits_pointsFinished = T43;
  assign T43 = outputReg_0_pointsFinished & T34;
  assign T44 = T27 ? T45 : outputReg_0_pointsFinished;
  assign T45 = inputReg_0_pointsFinished & T5;
  assign T46 = T50 && T47;
  assign T47 = T48;
  assign T48 = T49[1'h0/* 0*/:1'h0/* 0*/];
  assign T49 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T50 = T51 && io_in_valid;
  assign T51 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T52 = T46 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign io_out_bits_centeroidsFinished = T53;
  assign T53 = outputReg_0_centeroidsFinished & T34;
  assign T54 = T27 ? T55 : outputReg_0_centeroidsFinished;
  assign T55 = inputReg_0_centeroidsFinished & T5;
  assign T56 = T46 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T57 = T59 && T58;
  assign T58 = T40 == 8'hff/* 255*/;
  assign T59 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T60 = T104 ? 8'hff/* 255*/ : T61;
  assign T61 = T33 ? T64 : T62;
  assign T62 = T46 ? T63 : State_0;
  assign T63 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T64 = EmitReturnState_0 & T65;
  assign T65 = {4'h8/* 8*/{T34}};
  assign T66 = T93 || T67;
  assign T67 = T68 && T5;
  assign T68 = T20 && T69;
  assign T69 = ! T70;
  assign T70 = T71 >= 33'h9/* 9*/;
  assign T71 = {1'h0/* 0*/, T72};
  assign T72 = broadcastIndex_0 & T73;
  assign T73 = {6'h20/* 32*/{T5}};
  assign T74 = T75 || T67;
  assign T75 = T78 || T76;
  assign T76 = T77 && T5;
  assign T77 = T20 && T70;
  assign T78 = T46 || T79;
  assign T79 = T80 && T5;
  assign T80 = T28 && T81;
  assign T81 = mode == 32'h0/* 0*/;
  assign T82 = T84 || T83;
  assign T83 = T28 && T45;
  assign T84 = T28 && T55;
  assign T85 = T83 ? 32'h0/* 0*/ : T86;
  assign T86 = T84 ? 32'h1/* 1*/ : mode;
  assign T87 = T67 ? T92 : T88;
  assign T88 = T76 ? 32'h0/* 0*/ : T89;
  assign T89 = T79 ? T91 : T90;
  assign T90 = T46 ? 32'h0/* 0*/ : broadcastIndex_0;
  assign T91 = T72 + 32'h1/* 1*/;
  assign T92 = T72 + 32'h1/* 1*/;
  assign T93 = T94 || T76;
  assign T94 = T79 || T95;
  assign T95 = T96 && T5;
  assign T96 = T28 && T97;
  assign T97 = ! T81;
  assign T98 = T67 ? T103 : T99;
  assign T99 = T102 ? 8'h0/* 0*/ : T100;
  assign T100 = T79 ? T101 : EmitReturnState_0;
  assign T101 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T102 = T95 || T76;
  assign T103 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T104 = T27 || T4;
  assign T105 = subStateTh_0 == 1'h0/* 0*/;
  assign io_out_tag = T106;
  assign T106 = inputTag_0 & T107;
  assign T107 = {4'ha/* 10*/{T34}};
  assign T108 = T46 ? io_in_tag : inputTag_0;
  RREncode rThreadEncoder(
       .io_valid_0( T19 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_1 vThreadEncoder(
       .io_valid_0( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_2 sThreadEncoder(
       .io_valid_0( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_0 <= T60;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T10;
    if(T27) begin
      outputReg_0_pointsFinished <= T44;
    end
    if(T46) begin
      inputReg_0_pointsFinished <= T52;
    end
    if(T27) begin
      outputReg_0_centeroidsFinished <= T54;
    end
    if(T46) begin
      inputReg_0_centeroidsFinished <= T56;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T66) begin
      EmitReturnState_0 <= T98;
    end
    if(reset) begin
      broadcastIndex_0 <= 32'h0/* 0*/;
    end else if(T74) begin
      broadcastIndex_0 <= T87;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T82) begin
      mode <= T85;
    end
    if(T46) begin
      inputTag_0 <= T108;
    end
  end
endmodule

module RREncode_3(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_4(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_5(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire[31:0] T290;
  wire[31:0] T291;
  wire[31:0] T292;
  wire[31:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[31:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[31:0] T301;
  wire[31:0] T302;
  reg[31:0] centeroidIndex_1;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  wire[31:0] T322;
  wire[31:0] T323;
  wire[31:0] T324;
  wire[31:0] T325;
  reg[31:0] centeroidIndex_0;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  wire[31:0] T344;
  wire[31:0] T345;
  wire[31:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire[7:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire[7:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire[7:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire[7:0] T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire[7:0] T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire[7:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  reg[0:0] inputReg_2_pointsFinished;
  wire T400;
  wire T401;
  wire T402;
  reg[0:0] inputReg_1_pointsFinished;
  wire T403;
  wire T404;
  reg[0:0] inputReg_0_pointsFinished;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  reg[31:0] mode;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T421;
  wire T422;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T423;
  wire[31:0] T424;
  wire[31:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire[15:0] T438;
  wire[15:0] T439;
  wire[15:0] T440;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T441;
  wire[31:0] T442;
  wire[15:0] T443;
  wire[15:0] T444;
  wire[15:0] T445;
  reg[15:0] outputReg_1_centeroidIndex;
  wire[31:0] T446;
  wire[31:0] T447;
  wire[15:0] T448;
  wire[15:0] T449;
  reg[15:0] outputReg_0_centeroidIndex;
  wire[31:0] T450;
  wire[31:0] T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T347 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T300 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T289 && io_in_valid;
  assign T289 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T290 = T252 ? 32'h0/* 0*/ : T291;
  assign T291 = T259 ? T299 : T292;
  assign T292 = T261 ? 32'h0/* 0*/ : T293;
  assign T293 = T267 ? T298 : T294;
  assign T294 = T273 ? 32'h0/* 0*/ : T295;
  assign T295 = T279 ? T297 : T296;
  assign T296 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T297 = T248 + 32'h1/* 1*/;
  assign T298 = T248 + 32'h1/* 1*/;
  assign T299 = T248 + 32'h1/* 1*/;
  assign T300 = T324 | T301;
  assign T301 = centeroidIndex_1 & T302;
  assign T302 = {6'h20/* 32*/{T228}};
  assign T303 = T305 || T304;
  assign T304 = T253 && T228;
  assign T305 = T307 || T306;
  assign T306 = T254 && T228;
  assign T307 = T309 || T308;
  assign T308 = T262 && T228;
  assign T309 = T311 || T310;
  assign T310 = T268 && T228;
  assign T311 = T313 || T312;
  assign T312 = T274 && T228;
  assign T313 = T315 || T314;
  assign T314 = T280 && T228;
  assign T315 = T288 && T316;
  assign T316 = T286[1'h1/* 1*/];
  assign T317 = T304 ? 32'h0/* 0*/ : T318;
  assign T318 = T306 ? T299 : T319;
  assign T319 = T308 ? 32'h0/* 0*/ : T320;
  assign T320 = T310 ? T298 : T321;
  assign T321 = T312 ? 32'h0/* 0*/ : T322;
  assign T322 = T314 ? T297 : T323;
  assign T323 = T315 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T324 = centeroidIndex_0 & T325;
  assign T325 = {6'h20/* 32*/{T240}};
  assign T326 = T328 || T327;
  assign T327 = T253 && T240;
  assign T328 = T330 || T329;
  assign T329 = T254 && T240;
  assign T330 = T332 || T331;
  assign T331 = T262 && T240;
  assign T332 = T334 || T333;
  assign T333 = T268 && T240;
  assign T334 = T336 || T335;
  assign T335 = T274 && T240;
  assign T336 = T338 || T337;
  assign T337 = T280 && T240;
  assign T338 = T288 && T339;
  assign T339 = T286[1'h0/* 0*/];
  assign T340 = T327 ? 32'h0/* 0*/ : T341;
  assign T341 = T329 ? T299 : T342;
  assign T342 = T331 ? 32'h0/* 0*/ : T343;
  assign T343 = T333 ? T298 : T344;
  assign T344 = T335 ? 32'h0/* 0*/ : T345;
  assign T345 = T337 ? T297 : T346;
  assign T346 = T338 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T347 = T348 || T327;
  assign T348 = T349 || T331;
  assign T349 = T355 || T350;
  assign T350 = T351 && T240;
  assign T351 = T354 && T352;
  assign T352 = T232 == T353;
  assign T353 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T354 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T355 = T361 || T356;
  assign T356 = T357 && T240;
  assign T357 = T360 && T358;
  assign T358 = T232 == T359;
  assign T359 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T360 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T361 = T367 || T362;
  assign T362 = T363 && T240;
  assign T363 = T366 && T364;
  assign T364 = T232 == T365;
  assign T365 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T366 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T367 = T373 || T368;
  assign T368 = T369 && T240;
  assign T369 = T372 && T370;
  assign T370 = T232 == T371;
  assign T371 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T372 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T373 = T379 || T374;
  assign T374 = T375 && T240;
  assign T375 = T378 && T376;
  assign T376 = T232 == T377;
  assign T377 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T378 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T379 = T384 || T380;
  assign T380 = T381 && T240;
  assign T381 = T268 && T382;
  assign T382 = ! T383;
  assign T383 = T248 == 32'h5/* 5*/;
  assign T384 = T387 || T385;
  assign T385 = T386 && T240;
  assign T386 = T268 && T383;
  assign T387 = T393 || T388;
  assign T388 = T389 && T240;
  assign T389 = T392 && T390;
  assign T390 = T232 == T391;
  assign T391 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T392 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T393 = T394 || T335;
  assign T394 = T395 || T337;
  assign T395 = T410 || T396;
  assign T396 = T397 && T240;
  assign T397 = T406 && T398;
  assign T398 = T401 | T399;
  assign T399 = inputReg_2_pointsFinished & T5;
  assign T400 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T401 = T404 | T402;
  assign T402 = inputReg_1_pointsFinished & T228;
  assign T403 = T315 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T404 = inputReg_0_pointsFinished & T240;
  assign T405 = T338 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T426 || T411;
  assign T411 = T412 && T240;
  assign T412 = T406 && T413;
  assign T413 = mode == 32'h1/* 1*/;
  assign T414 = T415 || T397;
  assign T415 = T406 && T416;
  assign T416 = T419 | T417;
  assign T417 = inputReg_2_centeroidsFinished & T5;
  assign T418 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T419 = T422 | T420;
  assign T420 = inputReg_1_centeroidsFinished & T228;
  assign T421 = T315 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T422 = inputReg_0_centeroidsFinished & T240;
  assign T423 = T338 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T424 = T397 ? 32'h0/* 0*/ : T425;
  assign T425 = T415 ? 32'h1/* 1*/ : mode;
  assign T426 = T428 || T427;
  assign T427 = T415 && T240;
  assign T428 = T432 || T429;
  assign T429 = T430 && T240;
  assign T430 = T406 && T431;
  assign T431 = mode == 32'h0/* 0*/;
  assign T432 = T338 || T433;
  assign T433 = T434 && T97;
  assign T434 = T452 && io_out_ready;
  assign io_out_valid = T435;
  assign T435 = T437 && T436;
  assign T436 = T20 == 8'hff/* 255*/;
  assign T437 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T438;
  assign T438 = T443 | T439;
  assign T439 = outputReg_2_centeroidIndex & T440;
  assign T440 = {5'h10/* 16*/{T23}};
  assign T441 = T259 ? T248 : T442;
  assign T442 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T443 = T448 | T444;
  assign T444 = outputReg_1_centeroidIndex & T445;
  assign T445 = {5'h10/* 16*/{T87}};
  assign T446 = T306 ? T248 : T447;
  assign T447 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T448 = outputReg_0_centeroidIndex & T449;
  assign T449 = {5'h10/* 16*/{T97}};
  assign T450 = T329 ? T248 : T451;
  assign T451 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T327 ? 8'h0/* 0*/ : T458;
  assign T458 = T331 ? T501 : T459;
  assign T459 = T350 ? 8'h0/* 0*/ : T460;
  assign T460 = T356 ? T500 : T461;
  assign T461 = T362 ? T499 : T462;
  assign T462 = T368 ? T498 : T463;
  assign T463 = T374 ? T497 : T464;
  assign T464 = T380 ? T496 : T465;
  assign T465 = T385 ? T495 : T466;
  assign T466 = T388 ? T494 : T467;
  assign T467 = T335 ? T493 : T468;
  assign T468 = T337 ? 8'h0/* 0*/ : T469;
  assign T469 = T396 ? T492 : T470;
  assign T470 = T411 ? T491 : T471;
  assign T471 = T427 ? 8'h0/* 0*/ : T472;
  assign T472 = T429 ? T490 : T473;
  assign T473 = T433 ? T476 : T474;
  assign T474 = T338 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T304;
  assign T507 = T508 || T308;
  assign T508 = T510 || T509;
  assign T509 = T351 && T228;
  assign T510 = T512 || T511;
  assign T511 = T357 && T228;
  assign T512 = T514 || T513;
  assign T513 = T363 && T228;
  assign T514 = T516 || T515;
  assign T515 = T369 && T228;
  assign T516 = T518 || T517;
  assign T517 = T375 && T228;
  assign T518 = T520 || T519;
  assign T519 = T381 && T228;
  assign T520 = T522 || T521;
  assign T521 = T386 && T228;
  assign T522 = T524 || T523;
  assign T523 = T389 && T228;
  assign T524 = T525 || T312;
  assign T525 = T526 || T314;
  assign T526 = T528 || T527;
  assign T527 = T397 && T228;
  assign T528 = T530 || T529;
  assign T529 = T412 && T228;
  assign T530 = T532 || T531;
  assign T531 = T415 && T228;
  assign T532 = T534 || T533;
  assign T533 = T430 && T228;
  assign T534 = T315 || T535;
  assign T535 = T434 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T304 ? 8'h0/* 0*/ : T539;
  assign T539 = T308 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T312 ? T560 : T549;
  assign T549 = T314 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T315 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T351 && T5;
  assign T819 = T821 || T820;
  assign T820 = T357 && T5;
  assign T821 = T823 || T822;
  assign T822 = T363 && T5;
  assign T823 = T825 || T824;
  assign T824 = T369 && T5;
  assign T825 = T827 || T826;
  assign T826 = T375 && T5;
  assign T827 = T829 || T828;
  assign T828 = T381 && T5;
  assign T829 = T831 || T830;
  assign T830 = T386 && T5;
  assign T831 = T833 || T832;
  assign T832 = T389 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T397 && T5;
  assign T837 = T839 || T838;
  assign T838 = T412 && T5;
  assign T839 = T841 || T840;
  assign T840 = T415 && T5;
  assign T841 = T843 || T842;
  assign T842 = T430 && T5;
  assign T843 = T284 || T844;
  assign T844 = T434 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T315 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T338 ? io_in_tag : inputTag_0;
  RREncode_3 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_4 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_5 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T290;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T303) begin
      centeroidIndex_1 <= T317;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T326) begin
      centeroidIndex_0 <= T340;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T400;
    end
    if(T315) begin
      inputReg_1_pointsFinished <= T403;
    end
    if(T338) begin
      inputReg_0_pointsFinished <= T405;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T414) begin
      mode <= T424;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T418;
    end
    if(T315) begin
      inputReg_1_centeroidsFinished <= T421;
    end
    if(T338) begin
      inputReg_0_centeroidsFinished <= T423;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T441;
    end
    if(T306) begin
      outputReg_1_centeroidIndex <= T446;
    end
    if(T329) begin
      outputReg_0_centeroidIndex <= T450;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T315) begin
      inputTag_1 <= T894;
    end
    if(T338) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_6(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_7(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_8(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_6 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_7 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_8 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_1 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_2 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_2 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_3 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_2 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_3 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_4 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_3 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_5 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_4 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_5 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_6 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_5 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_6 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_7 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_6 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_7 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_8 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_7 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_8 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_8 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;
  assign T11 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_9 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_1(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_1 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_10 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_1 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_9 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  pcIn0_valid,
    input  pcIn0_bits_request,
    input [15:0] pcIn0_bits_moduleId,
    input [7:0] pcIn0_bits_portId,
    input [19:0] pcIn0_bits_pcValue,
    input [3:0] pcIn0_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_11 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_9 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_9(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_10(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_11(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_9 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_10 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_11 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_12(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_13(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_14(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_12 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_13 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_14 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_10 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_10 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_11 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_13 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_11 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_12 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_14 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_12 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_13 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_16(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_15 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_13 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_14 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_17(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_16 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_14 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_15 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_18(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_17 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_15 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_16(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_16(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_16 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_19(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_18 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_16 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_17(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_17(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_17 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_20(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_19 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_17 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_18(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_18(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_18 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_21(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_20 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_18 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_22(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_1 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_21 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_2(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_2 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_23(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_22 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_2 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_3(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_3 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_24(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_23 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_3 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_19(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_19(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_19 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_25(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_24 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_19 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_15(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_16(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_17(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_15 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_16 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_17 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_18(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_19(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_20(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_2(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_18 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_19 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_20 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_20(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_20(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_20 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_26(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_2 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_20 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_21(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_21(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_21 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_27(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_26 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_21 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_22(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_22(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_22 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_28(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_27 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_22 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_23(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_23(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_23 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_29(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_28 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_23 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_24(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_24(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_24 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_30(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_29 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_24 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_25(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_25(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_25 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_31(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_30 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_25 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_26(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_26(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_26 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_32(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_31 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_26 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_27(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_27(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_27 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_33(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_32 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_27 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_28(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_28(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_28 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_34(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_33 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_28 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_35(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_2 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_34 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_4(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_4 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_36(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_35 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_4 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_5(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_5 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_37(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_36 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_5 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_29(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_29(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_29 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_38(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_37 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_29 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_21(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_22(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_23(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_21 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_22 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_23 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_24(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_25(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_26(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_3(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_24 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_25 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_26 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_30(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_30(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_30 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_39(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_3 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_30 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_31(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_31(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_31 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_40(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_39 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_31 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_32(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_32(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_32 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_41(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_40 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_32 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_33(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_33(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_33 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_42(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_41 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_33 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_34(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_34(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_34 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_43(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_42 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_34 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_35(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_35(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_35 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_44(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_43 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_35 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_36(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_36(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_36 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_45(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_44 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_36 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_37(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_37(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_37 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_46(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_45 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_37 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_38(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_38(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_38 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_47(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_46 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_38 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_48(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_3 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_47 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_6(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_6 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_49(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_48 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_6 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_7(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_7 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_50(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_49 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_7 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_39(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_39(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_39 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_51(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_50 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_39 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_27(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_28(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_29(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_27 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_28 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_29 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_30(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_31(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_32(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_4(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_30 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_31 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_32 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_40(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_40(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_40 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_52(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_4 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_40 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_41(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_41(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_41 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_53(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_52 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_41 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_42(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_42(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_42 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_54(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_53 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_42 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_43(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_43(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_43 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_55(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_54 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_43 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_44(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_44(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_44 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_56(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_55 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_44 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_45(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_45(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_45 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_57(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_56 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_45 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_46(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_46(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_46 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_58(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_57 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_46 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_47(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_47(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_47 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_59(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_58 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_47 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_48(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_48(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_48 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_60(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_59 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_48 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_61(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_4 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_60 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_8(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_8 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_62(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_61 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_8 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_9(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_9 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_63(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_62 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_9 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_49(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_49(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_49 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_64(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_63 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_49 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_33(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_34(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_35(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_33 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_34 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_35 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_36(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_37(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_38(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_5(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_36 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_37 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_38 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_50(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_50(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_50 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_65(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_5 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_50 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_51(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_51(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_51 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_66(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_65 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_51 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_52(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_52(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_52 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_67(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_66 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_52 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_53(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_53(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_53 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_68(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_67 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_53 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_54(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_54(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_54 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_69(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_68 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_54 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_55(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_55(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_55 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_70(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_69 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_55 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_56(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_56(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_56 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_71(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_70 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_56 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_57(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_57(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_57 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_72(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_71 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_57 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_58(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_58(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_58 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_73(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_72 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_58 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_74(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_5 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_73 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_10(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_10(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_10 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_75(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_74 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_10 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_11(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_11(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_11 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_76(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_75 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_11 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_59(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_59(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_59 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_77(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_76 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_59 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_39(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_40(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_41(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_39 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_40 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_41 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_42(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_43(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_44(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_6(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_42 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_43 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_44 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_60(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_60(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_60 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_78(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_6 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_60 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_61(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_61(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_61 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_79(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_78 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_61 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_62(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_62(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_62 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_80(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_79 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_62 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_63(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_63(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_63 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_81(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_80 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_63 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_64(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_64(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_64 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_82(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_81 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_64 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_65(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_65(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_65 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_83(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_82 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_65 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_66(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_66(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_66 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_84(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_83 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_66 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_67(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_67(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_67 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_85(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_84 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_67 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_68(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_68(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_68 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_86(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_85 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_68 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_87(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_6 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_86 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_12(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_12(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_12 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_88(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_87 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_12 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_13(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_13(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_13 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_89(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_88 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_13 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_69(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_69(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_69 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_90(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_89 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_69 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_45(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_46(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_47(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_45 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_46 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_47 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_48(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_49(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_50(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_7(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_48 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_49 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_50 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_70(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_70(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_70 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_91(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_7 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_70 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_71(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_71(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_71 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_92(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_91 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_71 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_72(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_72(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_72 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_93(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_92 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_72 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_73(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_73(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_73 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_94(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_93 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_73 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_74(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_74(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_74 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_95(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_94 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_74 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_75(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_75(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_75 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_96(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_95 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_75 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_76(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_76(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_76 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_97(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_96 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_76 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_77(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_77(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_77 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_98(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_97 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_77 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_78(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_78(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_78 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_99(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_98 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_78 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_100(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_7 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_99 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_14(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_14(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_14 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_101(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_100 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_14 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_15(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_15(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_15 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_102(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_101 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_15 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_79(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_79(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_79 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_103(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_102 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_79 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_51(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_52(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_53(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_51 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_52 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_53 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_54(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_55(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_56(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_8(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_54 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_55 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_56 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_80(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_80(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_80 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_104(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_8 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_80 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_81(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_81(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_81 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_105(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_104 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_81 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_82(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_82(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_82 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_106(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_105 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_82 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_83(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_83(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_83 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_107(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_106 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_83 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_84(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_84(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_84 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_108(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_107 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_84 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_85(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_85(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_85 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_109(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_108 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_85 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_86(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_86(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_86 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_110(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_109 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_86 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_87(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_87(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_87 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_111(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_110 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_87 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_88(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_88(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_88 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_112(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_111 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_88 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_113(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_8 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_112 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_16(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_16(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_16 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_114(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_113 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_16 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_17(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_17(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_17 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_115(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_114 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_17 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_89(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_89(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_89 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_116(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_115 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_89 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_57(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_58(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module RREncode_59(input clk, input reset,
    input  io_valid_0,
    input  io_valid_1,
    input  io_valid_2,
    output[1:0] io_chosen,
    input  io_ready);

  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg[1:0] last_grant;
  wire T8;
  wire outValid;
  wire T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire[1:0] T14;

  assign io_chosen = choose;
  assign choose = T12 ? T11 : T0;
  assign T0 = T6 ? 2'h2/* 2*/ : T1;
  assign T1 = io_valid_0 ? T5 : T2;
  assign T2 = io_valid_1 ? T4 : T3;
  assign T3 = io_valid_2 ? 2'h2/* 2*/ : 2'h3/* 3*/;
  assign T4 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T5 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T6 = io_valid_2 && T7;
  assign T7 = 2'h2/* 2*/ > last_grant;
  assign T8 = outValid && io_ready;
  assign outValid = T9 || io_valid_2;
  assign T9 = io_valid_0 || io_valid_1;
  assign T10 = T8 ? choose : last_grant;
  assign T11 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T12 = io_valid_1 && T13;
  assign T13 = T14 > last_grant;
  assign T14 = {1'h0/* 0*/, 1'h1/* 1*/};

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0/* 0*/;
    end else if(T8) begin
      last_grant <= T10;
    end
  end
endmodule

module KEngine_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_distanceFU_req_ready,
    output mainOff_distanceFU_req_valid,
    output[63:0] mainOff_distanceFU_req_bits_in1_x,
    output[63:0] mainOff_distanceFU_req_bits_in1_y,
    output[63:0] mainOff_distanceFU_req_bits_in1_z,
    output[63:0] mainOff_distanceFU_req_bits_in2_x,
    output[63:0] mainOff_distanceFU_req_bits_in2_y,
    output[63:0] mainOff_distanceFU_req_bits_in2_z,
    output[9:0] mainOff_distanceFU_req_tag,
    output mainOff_distanceFU_rep_ready,
    input  mainOff_distanceFU_rep_valid,
    input [63:0] mainOff_distanceFU_rep_bits_out,
    input [9:0] mainOff_distanceFU_rep_tag,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire[1:0] sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_2;
  wire T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[5:0] T7;
  wire[1:0] vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_2;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_2;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire[7:0] T22;
  wire T23;
  wire[2:0] T24;
  wire[5:0] T25;
  wire[1:0] rThreadEncoder_io_chosen;
  wire T26;
  reg[0:0] subStateTh_2;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire AllOffloadsReady;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg[0:0] addPortHadReadyRequest;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg[0:0] add_ready_received;
  wire T45;
  wire T46;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire partialAccumulatorMemPort_req_valid;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[7:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[7:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  reg[0:0] partialAccumulatorMem_valid_received_2;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[9:0] T80;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T81;
  wire partialAccumulatorMemPort_rep_valid;
  wire T82;
  wire T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] partialAccumulatorMem_valid_received_1;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire[9:0] T92;
  wire T93;
  wire T94;
  wire[4:0] T95;
  wire T96;
  wire T97;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[9:0] T102;
  wire T103;
  wire T104;
  wire[4:0] T105;
  wire T106;
  wire T107;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T112;
  wire T113;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire centeroidMemPort_req_valid;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[7:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg[0:0] centeroidMem_valid_received_2;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire[9:0] T137;
  wire[9:0] centeroidMemPort_rep_tag;
  wire[9:0] centeroidMemPort_req_tag;
  wire[9:0] T138;
  wire centeroidMemPort_rep_valid;
  wire T139;
  wire T140;
  wire[4:0] T141;
  wire T142;
  wire T143;
  reg[0:0] centeroidMem_valid_received_1;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T148;
  wire T149;
  wire T150;
  wire[4:0] T151;
  wire T152;
  reg[0:0] centeroidMem_valid_received_0;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire[9:0] T157;
  wire T158;
  wire T159;
  wire[4:0] T160;
  wire T161;
  wire T162;
  reg[0:0] centeroidMemPortHadReadyRequest;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg[0:0] centeroidMem_ready_received;
  wire T167;
  wire T168;
  wire centeroidMemPort_req_ready;
  wire centeroidMemPort_rep_ready;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire distanceFUPort_req_valid;
  wire T173;
  wire T174;
  wire T175;
  wire[7:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] distanceFU_valid_received_2;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[9:0] distanceFUPort_rep_tag;
  wire distanceFUPort_rep_ready;
  wire[9:0] distanceFUPort_req_tag;
  wire[9:0] T187;
  wire distanceFUPort_rep_valid;
  wire T188;
  wire T189;
  wire[4:0] T190;
  wire T191;
  wire T192;
  reg[0:0] distanceFU_valid_received_1;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[9:0] T197;
  wire T198;
  wire T199;
  wire[4:0] T200;
  wire T201;
  reg[0:0] distanceFU_valid_received_0;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[9:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  reg[0:0] distanceFUPortHadReadyRequest;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg[0:0] distanceFU_ready_received;
  wire T216;
  wire T217;
  wire distanceFUPort_req_ready;
  wire T218;
  wire T219;
  reg[0:0] subStateTh_1;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire T225;
  reg[7:0] State_1;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[7:0] T237;
  wire[7:0] T238;
  wire[7:0] T239;
  wire T240;
  reg[7:0] State_0;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[31:0] T248;
  wire[31:0] T249;
  wire[31:0] T250;
  reg[31:0] centeroidIndex_2;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire[7:0] T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire[7:0] T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[7:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire[7:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire[2:0] T286;
  wire[5:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[15:0] T292;
  wire[15:0] T293;
  wire[15:0] T294;
  reg[15:0] outputReg_2_centeroidIndex;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[15:0] T297;
  wire[15:0] T298;
  wire[15:0] T299;
  reg[15:0] outputReg_1_centeroidIndex;
  wire T300;
  wire[31:0] T301;
  wire[31:0] T302;
  wire[15:0] T303;
  wire[15:0] T304;
  reg[15:0] outputReg_0_centeroidIndex;
  wire T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire T308;
  wire[31:0] T309;
  wire[31:0] T310;
  wire[31:0] T311;
  wire[31:0] T312;
  wire[31:0] T313;
  wire[31:0] T314;
  wire[31:0] T315;
  wire[31:0] T316;
  wire[31:0] T317;
  wire[31:0] T318;
  wire[31:0] T319;
  wire[31:0] T320;
  wire[31:0] T321;
  reg[31:0] centeroidIndex_1;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T340;
  wire[31:0] T341;
  wire[31:0] T342;
  wire[31:0] T343;
  reg[31:0] centeroidIndex_0;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire[31:0] T357;
  wire[31:0] T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire[31:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire[7:0] T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[7:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[7:0] T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[7:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[7:0] T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[7:0] T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] inputReg_2_pointsFinished;
  wire T417;
  wire T418;
  wire T419;
  reg[0:0] inputReg_1_pointsFinished;
  wire T420;
  wire T421;
  reg[0:0] inputReg_0_pointsFinished;
  wire T422;
  wire T423;
  wire T424;
  wire[7:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  reg[31:0] mode;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg[0:0] inputReg_2_centeroidsFinished;
  wire T435;
  wire T436;
  wire T437;
  reg[0:0] inputReg_1_centeroidsFinished;
  wire T438;
  wire T439;
  reg[0:0] inputReg_0_centeroidsFinished;
  wire T440;
  wire[31:0] T441;
  wire[31:0] T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire[7:0] T457;
  wire[7:0] T458;
  wire[7:0] T459;
  wire[7:0] T460;
  wire[7:0] T461;
  wire[7:0] T462;
  wire[7:0] T463;
  wire[7:0] T464;
  wire[7:0] T465;
  wire[7:0] T466;
  wire[7:0] T467;
  wire[7:0] T468;
  wire[7:0] T469;
  wire[7:0] T470;
  wire[7:0] T471;
  wire[7:0] T472;
  wire[7:0] T473;
  wire[7:0] T474;
  wire[7:0] T475;
  wire[7:0] T476;
  wire[7:0] T477;
  wire[7:0] T478;
  reg[7:0] EmitReturnState_2;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[7:0] T482;
  wire[7:0] T483;
  reg[7:0] EmitReturnState_1;
  wire[7:0] T484;
  wire[7:0] T485;
  wire[7:0] T486;
  wire[7:0] T487;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T488;
  wire[7:0] T489;
  wire[7:0] T490;
  wire[7:0] T491;
  wire[7:0] T492;
  wire[7:0] T493;
  wire[7:0] T494;
  wire[7:0] T495;
  wire[7:0] T496;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[7:0] T500;
  wire[7:0] T501;
  wire[7:0] T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[7:0] T536;
  wire[7:0] T537;
  wire[7:0] T538;
  wire[7:0] T539;
  wire[7:0] T540;
  wire[7:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  wire[7:0] T545;
  wire[7:0] T546;
  wire[7:0] T547;
  wire[7:0] T548;
  wire[7:0] T549;
  wire[7:0] T550;
  wire[7:0] T551;
  wire[7:0] T552;
  wire[7:0] T553;
  wire[7:0] T554;
  wire[7:0] T555;
  wire[7:0] T556;
  wire[7:0] T557;
  wire[7:0] T558;
  wire[7:0] T559;
  wire[7:0] T560;
  wire[7:0] T561;
  wire[7:0] T562;
  wire[7:0] T563;
  wire[7:0] T564;
  wire[7:0] T565;
  wire[7:0] T566;
  wire[7:0] T567;
  wire[7:0] T568;
  wire[7:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire T575;
  reg[0:0] subStateTh_0;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire[1:0] T586;
  wire T587;
  wire[7:0] T588;
  wire[7:0] T589;
  wire[7:0] T590;
  wire[7:0] T591;
  wire[7:0] T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[7:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[7:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  reg[0:0] add_valid_received_2;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire[9:0] T611;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T612;
  wire addPort_rep_valid;
  wire T613;
  wire T614;
  wire[4:0] T615;
  wire T616;
  wire T617;
  reg[0:0] add_valid_received_1;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[9:0] T622;
  wire T623;
  wire T624;
  wire[4:0] T625;
  wire T626;
  reg[0:0] add_valid_received_0;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire[4:0] T634;
  wire T635;
  wire T636;
  wire[4:0] T637;
  wire T638;
  wire T639;
  wire[4:0] T640;
  wire T641;
  wire T642;
  wire T643;
  wire[9:0] T644;
  wire T645;
  wire T646;
  wire T647;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_2;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[4:0] T652;
  wire T653;
  wire T654;
  wire[4:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[9:0] T659;
  wire T660;
  wire T661;
  wire T662;
  reg[0:0] centeroidMemPortHadValidRequest_2;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire[4:0] T667;
  wire T668;
  wire T669;
  wire[4:0] T670;
  wire T671;
  wire T672;
  wire T673;
  wire[9:0] T674;
  wire T675;
  wire T676;
  reg[0:0] distanceFUPortHadValidRequest_2;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire[4:0] T681;
  wire T682;
  wire T683;
  wire[4:0] T684;
  wire T685;
  wire T686;
  wire T687;
  wire[9:0] T688;
  wire T689;
  wire T690;
  wire AllOffloadsValid_1;
  wire T691;
  wire T692;
  wire T693;
  reg[0:0] addPortHadValidRequest_1;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire[4:0] T698;
  wire T699;
  wire T700;
  wire[4:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[9:0] T705;
  wire T706;
  wire T707;
  wire T708;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_1;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire[4:0] T713;
  wire T714;
  wire T715;
  wire[4:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire[9:0] T720;
  wire T721;
  wire T722;
  wire T723;
  reg[0:0] centeroidMemPortHadValidRequest_1;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[4:0] T728;
  wire T729;
  wire T730;
  wire[4:0] T731;
  wire T732;
  wire T733;
  wire T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  reg[0:0] distanceFUPortHadValidRequest_1;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[4:0] T742;
  wire T743;
  wire T744;
  wire[4:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire AllOffloadsValid_0;
  wire T752;
  wire T753;
  wire T754;
  reg[0:0] addPortHadValidRequest_0;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[4:0] T759;
  wire T760;
  wire T761;
  wire[4:0] T762;
  wire T763;
  wire T764;
  wire T765;
  wire[9:0] T766;
  wire T767;
  wire T768;
  wire T769;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[4:0] T774;
  wire T775;
  wire T776;
  wire[4:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  reg[0:0] centeroidMemPortHadValidRequest_0;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire[4:0] T789;
  wire T790;
  wire T791;
  wire[4:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[9:0] T796;
  wire T797;
  wire T798;
  reg[0:0] distanceFUPortHadValidRequest_0;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire[4:0] T803;
  wire T804;
  wire T805;
  wire[4:0] T806;
  wire T807;
  wire T808;
  wire T809;
  wire[9:0] T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire[7:0] T845;
  wire[7:0] T846;
  wire[7:0] T847;
  wire[7:0] T848;
  wire[7:0] T849;
  wire[7:0] T850;
  wire[7:0] T851;
  wire[7:0] T852;
  wire[7:0] T853;
  wire[7:0] T854;
  wire[7:0] T855;
  wire[7:0] T856;
  wire[7:0] T857;
  wire[7:0] T858;
  wire[7:0] T859;
  wire[7:0] T860;
  wire[7:0] T861;
  wire[7:0] T862;
  wire[7:0] T863;
  wire[7:0] T864;
  wire[7:0] T865;
  wire[7:0] T866;
  wire[7:0] T867;
  wire[7:0] T868;
  wire[7:0] T869;
  wire[7:0] T870;
  wire[7:0] T871;
  wire[7:0] T872;
  wire[7:0] T873;
  wire[7:0] T874;
  wire[7:0] T875;
  wire[7:0] T876;
  wire[7:0] T877;
  wire[7:0] T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire[9:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  reg[9:0] inputTag_2;
  wire[9:0] T890;
  wire[9:0] T891;
  wire[9:0] T892;
  wire[9:0] T893;
  reg[9:0] inputTag_1;
  wire[9:0] T894;
  wire[9:0] T895;
  wire[9:0] T896;
  reg[9:0] inputTag_0;
  wire[9:0] T897;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T1 = T879 && T2;
  assign T2 = State_2 == 8'h0/* 0*/;
  assign T3 = T813 || T4;
  assign T4 = T229 && T5;
  assign T5 = T6[2'h2/* 2*/];
  assign T6 = T7[2'h2/* 2*/:1'h0/* 0*/];
  assign T7 = 3'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T689 && AllOffloadsValid_2;
  assign AllOffloadsValid_2 = T9;
  assign T9 = T645 && T10;
  assign T10 = T641 || T11;
  assign T11 = ! addPortHadValidRequest_2;
  assign T12 = T638 && T13;
  assign T13 = addPortHadValidRequest_2 || T14;
  assign T14 = T636 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T603 && T16;
  assign T16 = T594 || T17;
  assign T17 = T593 && T18;
  assign T18 = T20 == T19;
  assign T19 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T20 = T588 | T21;
  assign T21 = State_2 & T22;
  assign T22 = {4'h8/* 8*/{T23}};
  assign T23 = T24[2'h2/* 2*/];
  assign T24 = T25[2'h2/* 2*/:1'h0/* 0*/];
  assign T25 = 3'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T26 = subStateTh_2 == 1'h0/* 0*/;
  assign T27 = T30 ? 1'h1/* 1*/ : T28;
  assign T28 = T29 ? 1'h0/* 0*/ : subStateTh_2;
  assign T29 = 2'h2/* 2*/ == vThreadEncoder_io_chosen;
  assign T30 = T32 && T31;
  assign T31 = State_2 != 8'hff/* 255*/;
  assign T32 = T34 && T33;
  assign T33 = State_2 != 8'h0/* 0*/;
  assign T34 = AllOffloadsReady && T35;
  assign T35 = 2'h2/* 2*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T36;
  assign T36 = T48 && T37;
  assign T37 = T44 || T38;
  assign T38 = T40 && T39;
  assign T39 = ! addPort_req_valid;
  assign T40 = ! addPortHadReadyRequest;
  assign T41 = T43 && T42;
  assign T42 = addPortHadReadyRequest || addPort_req_valid;
  assign T43 = ! AllOffloadsReady;
  assign T44 = addPort_req_ready || add_ready_received;
  assign T45 = T47 && T46;
  assign T46 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T47 = ! AllOffloadsReady;
  assign T48 = T115 && T49;
  assign T49 = T111 || T50;
  assign T50 = T107 && T51;
  assign T51 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T52;
  assign T52 = T72 && T53;
  assign T53 = T58 || T54;
  assign T54 = T57 && T55;
  assign T55 = T20 == T56;
  assign T56 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T57 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T58 = T63 || T59;
  assign T59 = T62 && T60;
  assign T60 = T20 == T61;
  assign T61 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T62 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T63 = T68 || T64;
  assign T64 = T67 && T65;
  assign T65 = T20 == T66;
  assign T66 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T67 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T68 = T71 && T69;
  assign T69 = T20 == T70;
  assign T70 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T72 = T106 && T73;
  assign T73 = ! T74;
  assign T74 = T85 | T75;
  assign T75 = partialAccumulatorMem_valid_received_2 & T23;
  assign T76 = T82 && T77;
  assign T77 = partialAccumulatorMem_valid_received_2 || T78;
  assign T78 = partialAccumulatorMemPort_rep_valid && T79;
  assign T79 = partialAccumulatorMemPort_rep_tag == T80;
  assign T80 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T81;
  assign T81 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T82 = ! T83;
  assign T83 = T84 == 5'h2/* 2*/;
  assign T84 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T85 = T96 | T86;
  assign T86 = partialAccumulatorMem_valid_received_1 & T87;
  assign T87 = T24[1'h1/* 1*/];
  assign T88 = T93 && T89;
  assign T89 = partialAccumulatorMem_valid_received_1 || T90;
  assign T90 = partialAccumulatorMemPort_rep_valid && T91;
  assign T91 = partialAccumulatorMemPort_rep_tag == T92;
  assign T92 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T93 = ! T94;
  assign T94 = T95 == 5'h1/* 1*/;
  assign T95 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T96 = partialAccumulatorMem_valid_received_0 & T97;
  assign T97 = T24[1'h0/* 0*/];
  assign T98 = T103 && T99;
  assign T99 = partialAccumulatorMem_valid_received_0 || T100;
  assign T100 = partialAccumulatorMemPort_rep_valid && T101;
  assign T101 = partialAccumulatorMemPort_rep_tag == T102;
  assign T102 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T103 = ! T104;
  assign T104 = T105 == 5'h0/* 0*/;
  assign T105 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T106 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T107 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T108 = T110 && T109;
  assign T109 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T110 = ! AllOffloadsReady;
  assign T111 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T112 = T114 && T113;
  assign T113 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T114 = ! AllOffloadsReady;
  assign T115 = T170 && T116;
  assign T116 = T166 || T117;
  assign T117 = T162 && T118;
  assign T118 = ! centeroidMemPort_req_valid;
  assign centeroidMemPort_req_valid = T119;
  assign T119 = T129 && T120;
  assign T120 = T125 || T121;
  assign T121 = T124 && T122;
  assign T122 = T20 == T123;
  assign T123 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T124 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T129 = T161 && T130;
  assign T130 = ! T131;
  assign T131 = T142 | T132;
  assign T132 = centeroidMem_valid_received_2 & T23;
  assign T133 = T139 && T134;
  assign T134 = centeroidMem_valid_received_2 || T135;
  assign T135 = centeroidMemPort_rep_valid && T136;
  assign T136 = centeroidMemPort_rep_tag == T137;
  assign T137 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign centeroidMemPort_rep_tag = mainOff_centeroidMem_rep_tag;
  assign mainOff_centeroidMem_req_tag = centeroidMemPort_req_tag;
  assign centeroidMemPort_req_tag = T138;
  assign T138 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign centeroidMemPort_rep_valid = mainOff_centeroidMem_rep_valid;
  assign mainOff_centeroidMem_req_valid = centeroidMemPort_req_valid;
  assign T139 = ! T140;
  assign T140 = T141 == 5'h2/* 2*/;
  assign T141 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T142 = T152 | T143;
  assign T143 = centeroidMem_valid_received_1 & T87;
  assign T144 = T149 && T145;
  assign T145 = centeroidMem_valid_received_1 || T146;
  assign T146 = centeroidMemPort_rep_valid && T147;
  assign T147 = centeroidMemPort_rep_tag == T148;
  assign T148 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T149 = ! T150;
  assign T150 = T151 == 5'h1/* 1*/;
  assign T151 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T152 = centeroidMem_valid_received_0 & T97;
  assign T153 = T158 && T154;
  assign T154 = centeroidMem_valid_received_0 || T155;
  assign T155 = centeroidMemPort_rep_valid && T156;
  assign T156 = centeroidMemPort_rep_tag == T157;
  assign T157 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T158 = ! T159;
  assign T159 = T160 == 5'h0/* 0*/;
  assign T160 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T161 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T162 = ! centeroidMemPortHadReadyRequest;
  assign T163 = T165 && T164;
  assign T164 = centeroidMemPortHadReadyRequest || centeroidMemPort_req_valid;
  assign T165 = ! AllOffloadsReady;
  assign T166 = centeroidMemPort_req_ready || centeroidMem_ready_received;
  assign T167 = T169 && T168;
  assign T168 = centeroidMem_ready_received || centeroidMemPort_req_ready;
  assign centeroidMemPort_req_ready = mainOff_centeroidMem_req_ready;
  assign mainOff_centeroidMem_rep_ready = centeroidMemPort_rep_ready;
  assign centeroidMemPort_rep_ready = 1'h1/* 1*/;
  assign T169 = ! AllOffloadsReady;
  assign T170 = T215 || T171;
  assign T171 = T211 && T172;
  assign T172 = ! distanceFUPort_req_valid;
  assign distanceFUPort_req_valid = T173;
  assign T173 = T178 && T174;
  assign T174 = T177 && T175;
  assign T175 = T20 == T176;
  assign T176 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T177 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T178 = T210 && T179;
  assign T179 = ! T180;
  assign T180 = T191 | T181;
  assign T181 = distanceFU_valid_received_2 & T23;
  assign T182 = T188 && T183;
  assign T183 = distanceFU_valid_received_2 || T184;
  assign T184 = distanceFUPort_rep_valid && T185;
  assign T185 = distanceFUPort_rep_tag == T186;
  assign T186 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign distanceFUPort_rep_tag = mainOff_distanceFU_rep_tag;
  assign mainOff_distanceFU_rep_ready = distanceFUPort_rep_ready;
  assign distanceFUPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_distanceFU_req_valid = distanceFUPort_req_valid;
  assign mainOff_distanceFU_req_tag = distanceFUPort_req_tag;
  assign distanceFUPort_req_tag = T187;
  assign T187 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign distanceFUPort_rep_valid = mainOff_distanceFU_rep_valid;
  assign T188 = ! T189;
  assign T189 = T190 == 5'h2/* 2*/;
  assign T190 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T191 = T201 | T192;
  assign T192 = distanceFU_valid_received_1 & T87;
  assign T193 = T198 && T194;
  assign T194 = distanceFU_valid_received_1 || T195;
  assign T195 = distanceFUPort_rep_valid && T196;
  assign T196 = distanceFUPort_rep_tag == T197;
  assign T197 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T198 = ! T199;
  assign T199 = T200 == 5'h1/* 1*/;
  assign T200 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T201 = distanceFU_valid_received_0 & T97;
  assign T202 = T207 && T203;
  assign T203 = distanceFU_valid_received_0 || T204;
  assign T204 = distanceFUPort_rep_valid && T205;
  assign T205 = distanceFUPort_rep_tag == T206;
  assign T206 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T207 = ! T208;
  assign T208 = T209 == 5'h0/* 0*/;
  assign T209 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T210 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T211 = ! distanceFUPortHadReadyRequest;
  assign T212 = T214 && T213;
  assign T213 = distanceFUPortHadReadyRequest || distanceFUPort_req_valid;
  assign T214 = ! AllOffloadsReady;
  assign T215 = distanceFUPort_req_ready || distanceFU_ready_received;
  assign T216 = T218 && T217;
  assign T217 = distanceFU_ready_received || distanceFUPort_req_ready;
  assign distanceFUPort_req_ready = mainOff_distanceFU_req_ready;
  assign T218 = ! AllOffloadsReady;
  assign T219 = subStateTh_1 == 1'h0/* 0*/;
  assign T220 = T224 ? 1'h1/* 1*/ : T221;
  assign T221 = T222 ? 1'h0/* 0*/ : subStateTh_1;
  assign T222 = T223 == vThreadEncoder_io_chosen;
  assign T223 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T224 = T570 && T225;
  assign T225 = State_1 != 8'hff/* 255*/;
  assign T226 = T504 || T227;
  assign T227 = T229 && T228;
  assign T228 = T6[1'h1/* 1*/];
  assign T229 = T503 && T230;
  assign T230 = T232 == T231;
  assign T231 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T232 = T235 | T233;
  assign T233 = State_2 & T234;
  assign T234 = {4'h8/* 8*/{T5}};
  assign T235 = T238 | T236;
  assign T236 = State_1 & T237;
  assign T237 = {4'h8/* 8*/{T228}};
  assign T238 = State_0 & T239;
  assign T239 = {4'h8/* 8*/{T240}};
  assign T240 = T6[1'h0/* 0*/];
  assign T241 = T243 || T242;
  assign T242 = T229 && T240;
  assign T243 = T364 || T244;
  assign T244 = T245 && T240;
  assign T245 = T254 && T246;
  assign T246 = ! T247;
  assign T247 = T248 == 32'h5/* 5*/;
  assign T248 = T319 | T249;
  assign T249 = centeroidIndex_2 & T250;
  assign T250 = {6'h20/* 32*/{T5}};
  assign T251 = T258 || T252;
  assign T252 = T253 && T5;
  assign T253 = T254 && T247;
  assign T254 = T257 && T255;
  assign T255 = T232 == T256;
  assign T256 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T257 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T258 = T260 || T259;
  assign T259 = T254 && T5;
  assign T260 = T266 || T261;
  assign T261 = T262 && T5;
  assign T262 = T265 && T263;
  assign T263 = T232 == T264;
  assign T264 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T265 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T266 = T272 || T267;
  assign T267 = T268 && T5;
  assign T268 = T271 && T269;
  assign T269 = T232 == T270;
  assign T270 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T271 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T272 = T278 || T273;
  assign T273 = T274 && T5;
  assign T274 = T277 && T275;
  assign T275 = T232 == T276;
  assign T276 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T277 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T278 = T284 || T279;
  assign T279 = T280 && T5;
  assign T280 = T283 && T281;
  assign T281 = T232 == T282;
  assign T282 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T283 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T284 = T288 && T285;
  assign T285 = T286[2'h2/* 2*/];
  assign T286 = T287[2'h2/* 2*/:1'h0/* 0*/];
  assign T287 = 3'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T288 = T308 && io_in_valid;
  assign io_out_valid = T289;
  assign T289 = T291 && T290;
  assign T290 = T20 == 8'hff/* 255*/;
  assign T291 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_bits_centeroidIndex = T292;
  assign T292 = T297 | T293;
  assign T293 = outputReg_2_centeroidIndex & T294;
  assign T294 = {5'h10/* 16*/{T23}};
  assign T295 = T259 ? T248 : T296;
  assign T296 = {16'h0/* 0*/, outputReg_2_centeroidIndex};
  assign T297 = T303 | T298;
  assign T298 = outputReg_1_centeroidIndex & T299;
  assign T299 = {5'h10/* 16*/{T87}};
  assign T300 = T254 && T228;
  assign T301 = T300 ? T248 : T302;
  assign T302 = {16'h0/* 0*/, outputReg_1_centeroidIndex};
  assign T303 = outputReg_0_centeroidIndex & T304;
  assign T304 = {5'h10/* 16*/{T97}};
  assign T305 = T254 && T240;
  assign T306 = T305 ? T248 : T307;
  assign T307 = {16'h0/* 0*/, outputReg_0_centeroidIndex};
  assign T308 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T309 = T252 ? 32'h0/* 0*/ : T310;
  assign T310 = T259 ? T318 : T311;
  assign T311 = T261 ? 32'h0/* 0*/ : T312;
  assign T312 = T267 ? T317 : T313;
  assign T313 = T273 ? 32'h0/* 0*/ : T314;
  assign T314 = T279 ? T316 : T315;
  assign T315 = T284 ? 32'h0/* 0*/ : centeroidIndex_2;
  assign T316 = T248 + 32'h1/* 1*/;
  assign T317 = T248 + 32'h1/* 1*/;
  assign T318 = T248 + 32'h1/* 1*/;
  assign T319 = T342 | T320;
  assign T320 = centeroidIndex_1 & T321;
  assign T321 = {6'h20/* 32*/{T228}};
  assign T322 = T324 || T323;
  assign T323 = T253 && T228;
  assign T324 = T325 || T300;
  assign T325 = T327 || T326;
  assign T326 = T262 && T228;
  assign T327 = T329 || T328;
  assign T328 = T268 && T228;
  assign T329 = T331 || T330;
  assign T330 = T274 && T228;
  assign T331 = T333 || T332;
  assign T332 = T280 && T228;
  assign T333 = T288 && T334;
  assign T334 = T286[1'h1/* 1*/];
  assign T335 = T323 ? 32'h0/* 0*/ : T336;
  assign T336 = T300 ? T318 : T337;
  assign T337 = T326 ? 32'h0/* 0*/ : T338;
  assign T338 = T328 ? T317 : T339;
  assign T339 = T330 ? 32'h0/* 0*/ : T340;
  assign T340 = T332 ? T316 : T341;
  assign T341 = T333 ? 32'h0/* 0*/ : centeroidIndex_1;
  assign T342 = centeroidIndex_0 & T343;
  assign T343 = {6'h20/* 32*/{T240}};
  assign T344 = T346 || T345;
  assign T345 = T253 && T240;
  assign T346 = T347 || T305;
  assign T347 = T349 || T348;
  assign T348 = T262 && T240;
  assign T349 = T351 || T350;
  assign T350 = T268 && T240;
  assign T351 = T353 || T352;
  assign T352 = T274 && T240;
  assign T353 = T355 || T354;
  assign T354 = T280 && T240;
  assign T355 = T288 && T356;
  assign T356 = T286[1'h0/* 0*/];
  assign T357 = T345 ? 32'h0/* 0*/ : T358;
  assign T358 = T305 ? T318 : T359;
  assign T359 = T348 ? 32'h0/* 0*/ : T360;
  assign T360 = T350 ? T317 : T361;
  assign T361 = T352 ? 32'h0/* 0*/ : T362;
  assign T362 = T354 ? T316 : T363;
  assign T363 = T355 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T364 = T365 || T345;
  assign T365 = T366 || T348;
  assign T366 = T372 || T367;
  assign T367 = T368 && T240;
  assign T368 = T371 && T369;
  assign T369 = T232 == T370;
  assign T370 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T371 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T372 = T378 || T373;
  assign T373 = T374 && T240;
  assign T374 = T377 && T375;
  assign T375 = T232 == T376;
  assign T376 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T377 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T378 = T384 || T379;
  assign T379 = T380 && T240;
  assign T380 = T383 && T381;
  assign T381 = T232 == T382;
  assign T382 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T383 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T384 = T390 || T385;
  assign T385 = T386 && T240;
  assign T386 = T389 && T387;
  assign T387 = T232 == T388;
  assign T388 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T389 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T390 = T396 || T391;
  assign T391 = T392 && T240;
  assign T392 = T395 && T393;
  assign T393 = T232 == T394;
  assign T394 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T395 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T396 = T401 || T397;
  assign T397 = T398 && T240;
  assign T398 = T268 && T399;
  assign T399 = ! T400;
  assign T400 = T248 == 32'h5/* 5*/;
  assign T401 = T404 || T402;
  assign T402 = T403 && T240;
  assign T403 = T268 && T400;
  assign T404 = T410 || T405;
  assign T405 = T406 && T240;
  assign T406 = T409 && T407;
  assign T407 = T232 == T408;
  assign T408 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T409 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T410 = T411 || T352;
  assign T411 = T412 || T354;
  assign T412 = T427 || T413;
  assign T413 = T414 && T240;
  assign T414 = T423 && T415;
  assign T415 = T418 | T416;
  assign T416 = inputReg_2_pointsFinished & T5;
  assign T417 = T284 ? io_in_bits_pointsFinished : inputReg_2_pointsFinished;
  assign T418 = T421 | T419;
  assign T419 = inputReg_1_pointsFinished & T228;
  assign T420 = T333 ? io_in_bits_pointsFinished : inputReg_1_pointsFinished;
  assign T421 = inputReg_0_pointsFinished & T240;
  assign T422 = T355 ? io_in_bits_pointsFinished : inputReg_0_pointsFinished;
  assign T423 = T426 && T424;
  assign T424 = T232 == T425;
  assign T425 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T426 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T427 = T443 || T428;
  assign T428 = T429 && T240;
  assign T429 = T423 && T430;
  assign T430 = mode == 32'h1/* 1*/;
  assign T431 = T432 || T414;
  assign T432 = T423 && T433;
  assign T433 = T436 | T434;
  assign T434 = inputReg_2_centeroidsFinished & T5;
  assign T435 = T284 ? io_in_bits_centeroidsFinished : inputReg_2_centeroidsFinished;
  assign T436 = T439 | T437;
  assign T437 = inputReg_1_centeroidsFinished & T228;
  assign T438 = T333 ? io_in_bits_centeroidsFinished : inputReg_1_centeroidsFinished;
  assign T439 = inputReg_0_centeroidsFinished & T240;
  assign T440 = T355 ? io_in_bits_centeroidsFinished : inputReg_0_centeroidsFinished;
  assign T441 = T414 ? 32'h0/* 0*/ : T442;
  assign T442 = T432 ? 32'h1/* 1*/ : mode;
  assign T443 = T445 || T444;
  assign T444 = T432 && T240;
  assign T445 = T449 || T446;
  assign T446 = T447 && T240;
  assign T447 = T423 && T448;
  assign T448 = mode == 32'h0/* 0*/;
  assign T449 = T355 || T450;
  assign T450 = T451 && T97;
  assign T451 = T452 && io_out_ready;
  assign T452 = T454 && T453;
  assign T453 = T20 == 8'hff/* 255*/;
  assign T454 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T455 = T242 ? 8'hff/* 255*/ : T456;
  assign T456 = T244 ? T502 : T457;
  assign T457 = T345 ? 8'h0/* 0*/ : T458;
  assign T458 = T348 ? T501 : T459;
  assign T459 = T367 ? 8'h0/* 0*/ : T460;
  assign T460 = T373 ? T500 : T461;
  assign T461 = T379 ? T499 : T462;
  assign T462 = T385 ? T498 : T463;
  assign T463 = T391 ? T497 : T464;
  assign T464 = T397 ? T496 : T465;
  assign T465 = T402 ? T495 : T466;
  assign T466 = T405 ? T494 : T467;
  assign T467 = T352 ? T493 : T468;
  assign T468 = T354 ? 8'h0/* 0*/ : T469;
  assign T469 = T413 ? T492 : T470;
  assign T470 = T428 ? T491 : T471;
  assign T471 = T444 ? 8'h0/* 0*/ : T472;
  assign T472 = T446 ? T490 : T473;
  assign T473 = T450 ? T476 : T474;
  assign T474 = T355 ? T475 : State_0;
  assign T475 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T476 = T481 | T477;
  assign T477 = EmitReturnState_2 & T478;
  assign T478 = {4'h8/* 8*/{T23}};
  assign T479 = T4 ? T480 : EmitReturnState_2;
  assign T480 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T481 = T486 | T482;
  assign T482 = EmitReturnState_1 & T483;
  assign T483 = {4'h8/* 8*/{T87}};
  assign T484 = T227 ? T485 : EmitReturnState_1;
  assign T485 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T486 = EmitReturnState_0 & T487;
  assign T487 = {4'h8/* 8*/{T97}};
  assign T488 = T242 ? T489 : EmitReturnState_0;
  assign T489 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T490 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T491 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T492 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T493 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T494 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T495 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T496 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T497 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T498 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T499 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T500 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T501 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T502 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T503 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T504 = T506 || T505;
  assign T505 = T245 && T228;
  assign T506 = T507 || T323;
  assign T507 = T508 || T326;
  assign T508 = T510 || T509;
  assign T509 = T368 && T228;
  assign T510 = T512 || T511;
  assign T511 = T374 && T228;
  assign T512 = T514 || T513;
  assign T513 = T380 && T228;
  assign T514 = T516 || T515;
  assign T515 = T386 && T228;
  assign T516 = T518 || T517;
  assign T517 = T392 && T228;
  assign T518 = T520 || T519;
  assign T519 = T398 && T228;
  assign T520 = T522 || T521;
  assign T521 = T403 && T228;
  assign T522 = T524 || T523;
  assign T523 = T406 && T228;
  assign T524 = T525 || T330;
  assign T525 = T526 || T332;
  assign T526 = T528 || T527;
  assign T527 = T414 && T228;
  assign T528 = T530 || T529;
  assign T529 = T429 && T228;
  assign T530 = T532 || T531;
  assign T531 = T432 && T228;
  assign T532 = T534 || T533;
  assign T533 = T447 && T228;
  assign T534 = T333 || T535;
  assign T535 = T451 && T87;
  assign T536 = T227 ? 8'hff/* 255*/ : T537;
  assign T537 = T505 ? T569 : T538;
  assign T538 = T323 ? 8'h0/* 0*/ : T539;
  assign T539 = T326 ? T568 : T540;
  assign T540 = T509 ? 8'h0/* 0*/ : T541;
  assign T541 = T511 ? T567 : T542;
  assign T542 = T513 ? T566 : T543;
  assign T543 = T515 ? T565 : T544;
  assign T544 = T517 ? T564 : T545;
  assign T545 = T519 ? T563 : T546;
  assign T546 = T521 ? T562 : T547;
  assign T547 = T523 ? T561 : T548;
  assign T548 = T330 ? T560 : T549;
  assign T549 = T332 ? 8'h0/* 0*/ : T550;
  assign T550 = T527 ? T559 : T551;
  assign T551 = T529 ? T558 : T552;
  assign T552 = T531 ? 8'h0/* 0*/ : T553;
  assign T553 = T533 ? T557 : T554;
  assign T554 = T535 ? T476 : T555;
  assign T555 = T333 ? T556 : State_1;
  assign T556 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T557 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T558 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T559 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T560 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T561 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T562 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T563 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T564 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T565 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T566 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T567 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T568 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T569 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T570 = T572 && T571;
  assign T571 = State_1 != 8'h0/* 0*/;
  assign T572 = AllOffloadsReady && T573;
  assign T573 = T574 == rThreadEncoder_io_chosen;
  assign T574 = {1'h0/* 0*/, 1'h1/* 1*/};
  assign T575 = subStateTh_0 == 1'h0/* 0*/;
  assign T576 = T580 ? 1'h1/* 1*/ : T577;
  assign T577 = T578 ? 1'h0/* 0*/ : subStateTh_0;
  assign T578 = T579 == vThreadEncoder_io_chosen;
  assign T579 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T580 = T582 && T581;
  assign T581 = State_0 != 8'hff/* 255*/;
  assign T582 = T584 && T583;
  assign T583 = State_0 != 8'h0/* 0*/;
  assign T584 = AllOffloadsReady && T585;
  assign T585 = T586 == rThreadEncoder_io_chosen;
  assign T586 = {1'h0/* 0*/, 1'h0/* 0*/};
  assign T587 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T588 = T591 | T589;
  assign T589 = State_1 & T590;
  assign T590 = {4'h8/* 8*/{T87}};
  assign T591 = State_0 & T592;
  assign T592 = {4'h8/* 8*/{T97}};
  assign T593 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T594 = T599 || T595;
  assign T595 = T598 && T596;
  assign T596 = T20 == T597;
  assign T597 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T598 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T599 = T602 && T600;
  assign T600 = T20 == T601;
  assign T601 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T602 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T603 = T635 && T604;
  assign T604 = ! T605;
  assign T605 = T616 | T606;
  assign T606 = add_valid_received_2 & T23;
  assign T607 = T613 && T608;
  assign T608 = add_valid_received_2 || T609;
  assign T609 = addPort_rep_valid && T610;
  assign T610 = addPort_rep_tag == T611;
  assign T611 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T612;
  assign T612 = {8'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T613 = ! T614;
  assign T614 = T615 == 5'h2/* 2*/;
  assign T615 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T616 = T626 | T617;
  assign T617 = add_valid_received_1 & T87;
  assign T618 = T623 && T619;
  assign T619 = add_valid_received_1 || T620;
  assign T620 = addPort_rep_valid && T621;
  assign T621 = addPort_rep_tag == T622;
  assign T622 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T623 = ! T624;
  assign T624 = T625 == 5'h1/* 1*/;
  assign T625 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T626 = add_valid_received_0 & T97;
  assign T627 = T632 && T628;
  assign T628 = add_valid_received_0 || T629;
  assign T629 = addPort_rep_valid && T630;
  assign T630 = addPort_rep_tag == T631;
  assign T631 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T632 = ! T633;
  assign T633 = T634 == 5'h0/* 0*/;
  assign T634 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T635 = rThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T636 = 5'h2/* 2*/ == T637;
  assign T637 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T638 = ! T639;
  assign T639 = T640 == 5'h2/* 2*/;
  assign T640 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T641 = T642 || add_valid_received_2;
  assign T642 = addPort_rep_valid && T643;
  assign T643 = addPort_rep_tag == T644;
  assign T644 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T645 = T660 && T646;
  assign T646 = T656 || T647;
  assign T647 = ! partialAccumulatorMemPortHadValidRequest_2;
  assign T648 = T653 && T649;
  assign T649 = partialAccumulatorMemPortHadValidRequest_2 || T650;
  assign T650 = T651 && partialAccumulatorMemPort_req_valid;
  assign T651 = 5'h2/* 2*/ == T652;
  assign T652 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T653 = ! T654;
  assign T654 = T655 == 5'h2/* 2*/;
  assign T655 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T656 = T657 || partialAccumulatorMem_valid_received_2;
  assign T657 = partialAccumulatorMemPort_rep_valid && T658;
  assign T658 = partialAccumulatorMemPort_rep_tag == T659;
  assign T659 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T660 = T675 && T661;
  assign T661 = T671 || T662;
  assign T662 = ! centeroidMemPortHadValidRequest_2;
  assign T663 = T668 && T664;
  assign T664 = centeroidMemPortHadValidRequest_2 || T665;
  assign T665 = T666 && centeroidMemPort_req_valid;
  assign T666 = 5'h2/* 2*/ == T667;
  assign T667 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T668 = ! T669;
  assign T669 = T670 == 5'h2/* 2*/;
  assign T670 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T671 = T672 || centeroidMem_valid_received_2;
  assign T672 = centeroidMemPort_rep_valid && T673;
  assign T673 = centeroidMemPort_rep_tag == T674;
  assign T674 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T675 = T685 || T676;
  assign T676 = ! distanceFUPortHadValidRequest_2;
  assign T677 = T682 && T678;
  assign T678 = distanceFUPortHadValidRequest_2 || T679;
  assign T679 = T680 && distanceFUPort_req_valid;
  assign T680 = 5'h2/* 2*/ == T681;
  assign T681 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T682 = ! T683;
  assign T683 = T684 == 5'h2/* 2*/;
  assign T684 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T685 = T686 || distanceFU_valid_received_2;
  assign T686 = distanceFUPort_rep_valid && T687;
  assign T687 = distanceFUPort_rep_tag == T688;
  assign T688 = {5'h0/* 0*/, 5'h2/* 2*/};
  assign T689 = subStateTh_2 == 1'h1/* 1*/;
  assign T690 = T750 && AllOffloadsValid_1;
  assign AllOffloadsValid_1 = T691;
  assign T691 = T706 && T692;
  assign T692 = T702 || T693;
  assign T693 = ! addPortHadValidRequest_1;
  assign T694 = T699 && T695;
  assign T695 = addPortHadValidRequest_1 || T696;
  assign T696 = T697 && addPort_req_valid;
  assign T697 = 5'h1/* 1*/ == T698;
  assign T698 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T699 = ! T700;
  assign T700 = T701 == 5'h1/* 1*/;
  assign T701 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T702 = T703 || add_valid_received_1;
  assign T703 = addPort_rep_valid && T704;
  assign T704 = addPort_rep_tag == T705;
  assign T705 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T706 = T721 && T707;
  assign T707 = T717 || T708;
  assign T708 = ! partialAccumulatorMemPortHadValidRequest_1;
  assign T709 = T714 && T710;
  assign T710 = partialAccumulatorMemPortHadValidRequest_1 || T711;
  assign T711 = T712 && partialAccumulatorMemPort_req_valid;
  assign T712 = 5'h1/* 1*/ == T713;
  assign T713 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T714 = ! T715;
  assign T715 = T716 == 5'h1/* 1*/;
  assign T716 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T717 = T718 || partialAccumulatorMem_valid_received_1;
  assign T718 = partialAccumulatorMemPort_rep_valid && T719;
  assign T719 = partialAccumulatorMemPort_rep_tag == T720;
  assign T720 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T721 = T736 && T722;
  assign T722 = T732 || T723;
  assign T723 = ! centeroidMemPortHadValidRequest_1;
  assign T724 = T729 && T725;
  assign T725 = centeroidMemPortHadValidRequest_1 || T726;
  assign T726 = T727 && centeroidMemPort_req_valid;
  assign T727 = 5'h1/* 1*/ == T728;
  assign T728 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T729 = ! T730;
  assign T730 = T731 == 5'h1/* 1*/;
  assign T731 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T732 = T733 || centeroidMem_valid_received_1;
  assign T733 = centeroidMemPort_rep_valid && T734;
  assign T734 = centeroidMemPort_rep_tag == T735;
  assign T735 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T736 = T746 || T737;
  assign T737 = ! distanceFUPortHadValidRequest_1;
  assign T738 = T743 && T739;
  assign T739 = distanceFUPortHadValidRequest_1 || T740;
  assign T740 = T741 && distanceFUPort_req_valid;
  assign T741 = 5'h1/* 1*/ == T742;
  assign T742 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T743 = ! T744;
  assign T744 = T745 == 5'h1/* 1*/;
  assign T745 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T746 = T747 || distanceFU_valid_received_1;
  assign T747 = distanceFUPort_rep_valid && T748;
  assign T748 = distanceFUPort_rep_tag == T749;
  assign T749 = {5'h0/* 0*/, 5'h1/* 1*/};
  assign T750 = subStateTh_1 == 1'h1/* 1*/;
  assign T751 = T811 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T752;
  assign T752 = T767 && T753;
  assign T753 = T763 || T754;
  assign T754 = ! addPortHadValidRequest_0;
  assign T755 = T760 && T756;
  assign T756 = addPortHadValidRequest_0 || T757;
  assign T757 = T758 && addPort_req_valid;
  assign T758 = 5'h0/* 0*/ == T759;
  assign T759 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T760 = ! T761;
  assign T761 = T762 == 5'h0/* 0*/;
  assign T762 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T763 = T764 || add_valid_received_0;
  assign T764 = addPort_rep_valid && T765;
  assign T765 = addPort_rep_tag == T766;
  assign T766 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T767 = T782 && T768;
  assign T768 = T778 || T769;
  assign T769 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T770 = T775 && T771;
  assign T771 = partialAccumulatorMemPortHadValidRequest_0 || T772;
  assign T772 = T773 && partialAccumulatorMemPort_req_valid;
  assign T773 = 5'h0/* 0*/ == T774;
  assign T774 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T775 = ! T776;
  assign T776 = T777 == 5'h0/* 0*/;
  assign T777 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T778 = T779 || partialAccumulatorMem_valid_received_0;
  assign T779 = partialAccumulatorMemPort_rep_valid && T780;
  assign T780 = partialAccumulatorMemPort_rep_tag == T781;
  assign T781 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T782 = T797 && T783;
  assign T783 = T793 || T784;
  assign T784 = ! centeroidMemPortHadValidRequest_0;
  assign T785 = T790 && T786;
  assign T786 = centeroidMemPortHadValidRequest_0 || T787;
  assign T787 = T788 && centeroidMemPort_req_valid;
  assign T788 = 5'h0/* 0*/ == T789;
  assign T789 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T790 = ! T791;
  assign T791 = T792 == 5'h0/* 0*/;
  assign T792 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T793 = T794 || centeroidMem_valid_received_0;
  assign T794 = centeroidMemPort_rep_valid && T795;
  assign T795 = centeroidMemPort_rep_tag == T796;
  assign T796 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T797 = T807 || T798;
  assign T798 = ! distanceFUPortHadValidRequest_0;
  assign T799 = T804 && T800;
  assign T800 = distanceFUPortHadValidRequest_0 || T801;
  assign T801 = T802 && distanceFUPort_req_valid;
  assign T802 = 5'h0/* 0*/ == T803;
  assign T803 = {3'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T804 = ! T805;
  assign T805 = T806 == 5'h0/* 0*/;
  assign T806 = {3'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T807 = T808 || distanceFU_valid_received_0;
  assign T808 = distanceFUPort_rep_valid && T809;
  assign T809 = distanceFUPort_rep_tag == T810;
  assign T810 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T811 = subStateTh_0 == 1'h1/* 1*/;
  assign T812 = vThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign T813 = T815 || T814;
  assign T814 = T245 && T5;
  assign T815 = T816 || T252;
  assign T816 = T817 || T261;
  assign T817 = T819 || T818;
  assign T818 = T368 && T5;
  assign T819 = T821 || T820;
  assign T820 = T374 && T5;
  assign T821 = T823 || T822;
  assign T822 = T380 && T5;
  assign T823 = T825 || T824;
  assign T824 = T386 && T5;
  assign T825 = T827 || T826;
  assign T826 = T392 && T5;
  assign T827 = T829 || T828;
  assign T828 = T398 && T5;
  assign T829 = T831 || T830;
  assign T830 = T403 && T5;
  assign T831 = T833 || T832;
  assign T832 = T406 && T5;
  assign T833 = T834 || T273;
  assign T834 = T835 || T279;
  assign T835 = T837 || T836;
  assign T836 = T414 && T5;
  assign T837 = T839 || T838;
  assign T838 = T429 && T5;
  assign T839 = T841 || T840;
  assign T840 = T432 && T5;
  assign T841 = T843 || T842;
  assign T842 = T447 && T5;
  assign T843 = T284 || T844;
  assign T844 = T451 && T23;
  assign T845 = T4 ? 8'hff/* 255*/ : T846;
  assign T846 = T814 ? T878 : T847;
  assign T847 = T252 ? 8'h0/* 0*/ : T848;
  assign T848 = T261 ? T877 : T849;
  assign T849 = T818 ? 8'h0/* 0*/ : T850;
  assign T850 = T820 ? T876 : T851;
  assign T851 = T822 ? T875 : T852;
  assign T852 = T824 ? T874 : T853;
  assign T853 = T826 ? T873 : T854;
  assign T854 = T828 ? T872 : T855;
  assign T855 = T830 ? T871 : T856;
  assign T856 = T832 ? T870 : T857;
  assign T857 = T273 ? T869 : T858;
  assign T858 = T279 ? 8'h0/* 0*/ : T859;
  assign T859 = T836 ? T868 : T860;
  assign T860 = T838 ? T867 : T861;
  assign T861 = T840 ? 8'h0/* 0*/ : T862;
  assign T862 = T842 ? T866 : T863;
  assign T863 = T844 ? T476 : T864;
  assign T864 = T284 ? T865 : State_2;
  assign T865 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T866 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T867 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T868 = {4'h0/* 0*/, 4'hb/* 11*/};
  assign T869 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T870 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T871 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T872 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T873 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign T874 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign T875 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign T876 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign T877 = {4'h0/* 0*/, 4'hc/* 12*/};
  assign T878 = {4'h0/* 0*/, 4'hd/* 13*/};
  assign T879 = subStateTh_2 == 1'h0/* 0*/;
  assign T880 = T882 && T881;
  assign T881 = State_1 == 8'h0/* 0*/;
  assign T882 = subStateTh_1 == 1'h0/* 0*/;
  assign T883 = T885 && T884;
  assign T884 = State_0 == 8'h0/* 0*/;
  assign T885 = subStateTh_0 == 1'h0/* 0*/;
  assign T886 = sThreadEncoder_io_chosen != 2'h3/* 3*/;
  assign io_out_tag = T887;
  assign T887 = T891 | T888;
  assign T888 = inputTag_2 & T889;
  assign T889 = {4'ha/* 10*/{T23}};
  assign T890 = T284 ? io_in_tag : inputTag_2;
  assign T891 = T895 | T892;
  assign T892 = inputTag_1 & T893;
  assign T893 = {4'ha/* 10*/{T87}};
  assign T894 = T333 ? io_in_tag : inputTag_1;
  assign T895 = inputTag_0 & T896;
  assign T896 = {4'ha/* 10*/{T97}};
  assign T897 = T355 ? io_in_tag : inputTag_0;
  RREncode_57 rThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T575 ),
       .io_valid_1( T219 ),
       .io_valid_2( T26 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready( T587 ));
  RREncode_58 vThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T751 ),
       .io_valid_1( T690 ),
       .io_valid_2( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready( T812 ));
  RREncode_59 sThreadEncoder(.clk(clk), .reset(reset),
       .io_valid_0( T883 ),
       .io_valid_1( T880 ),
       .io_valid_2( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready( T886 ));

  always @(posedge clk) begin
    if(reset) begin
      State_2 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_2 <= T845;
    end
    addPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_2 <= reset ? 1'h0/* 0*/ : T27;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T41;
    add_ready_received <= reset ? 1'h0/* 0*/ : T45;
    partialAccumulatorMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T76;
    partialAccumulatorMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T88;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T98;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T108;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T112;
    centeroidMem_valid_received_2 <= reset ? 1'h0/* 0*/ : T133;
    centeroidMem_valid_received_1 <= reset ? 1'h0/* 0*/ : T144;
    centeroidMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T153;
    centeroidMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T163;
    centeroidMem_ready_received <= reset ? 1'h0/* 0*/ : T167;
    distanceFU_valid_received_2 <= reset ? 1'h0/* 0*/ : T182;
    distanceFU_valid_received_1 <= reset ? 1'h0/* 0*/ : T193;
    distanceFU_valid_received_0 <= reset ? 1'h0/* 0*/ : T202;
    distanceFUPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T212;
    distanceFU_ready_received <= reset ? 1'h0/* 0*/ : T216;
    subStateTh_1 <= reset ? 1'h0/* 0*/ : T220;
    if(reset) begin
      State_1 <= 8'h0/* 0*/;
    end else if(T226) begin
      State_1 <= T536;
    end
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T241) begin
      State_0 <= T455;
    end
    if(reset) begin
      centeroidIndex_2 <= 32'h0/* 0*/;
    end else if(T251) begin
      centeroidIndex_2 <= T309;
    end
    if(T259) begin
      outputReg_2_centeroidIndex <= T295;
    end
    if(T300) begin
      outputReg_1_centeroidIndex <= T301;
    end
    if(T305) begin
      outputReg_0_centeroidIndex <= T306;
    end
    if(reset) begin
      centeroidIndex_1 <= 32'h0/* 0*/;
    end else if(T322) begin
      centeroidIndex_1 <= T335;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T344) begin
      centeroidIndex_0 <= T357;
    end
    if(T284) begin
      inputReg_2_pointsFinished <= T417;
    end
    if(T333) begin
      inputReg_1_pointsFinished <= T420;
    end
    if(T355) begin
      inputReg_0_pointsFinished <= T422;
    end
    if(reset) begin
      mode <= 32'h0/* 0*/;
    end else if(T431) begin
      mode <= T441;
    end
    if(T284) begin
      inputReg_2_centeroidsFinished <= T435;
    end
    if(T333) begin
      inputReg_1_centeroidsFinished <= T438;
    end
    if(T355) begin
      inputReg_0_centeroidsFinished <= T440;
    end
    if(reset) begin
      EmitReturnState_2 <= 8'h0/* 0*/;
    end else if(T4) begin
      EmitReturnState_2 <= T479;
    end
    if(reset) begin
      EmitReturnState_1 <= 8'h0/* 0*/;
    end else if(T227) begin
      EmitReturnState_1 <= T484;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T242) begin
      EmitReturnState_0 <= T488;
    end
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T576;
    add_valid_received_2 <= reset ? 1'h0/* 0*/ : T607;
    add_valid_received_1 <= reset ? 1'h0/* 0*/ : T618;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T627;
    partialAccumulatorMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T648;
    centeroidMemPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T663;
    distanceFUPortHadValidRequest_2 <= reset ? 1'h0/* 0*/ : T677;
    addPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T694;
    partialAccumulatorMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T709;
    centeroidMemPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T724;
    distanceFUPortHadValidRequest_1 <= reset ? 1'h0/* 0*/ : T738;
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T755;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T770;
    centeroidMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T785;
    distanceFUPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T799;
    if(T284) begin
      inputTag_2 <= T890;
    end
    if(T333) begin
      inputTag_1 <= T894;
    end
    if(T355) begin
      inputTag_0 <= T897;
    end
  end
endmodule

module RREncode_60(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_61(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_62(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module distanceFU_9(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub1_req_ready,
    output mainOff_sub1_req_valid,
    output[63:0] mainOff_sub1_req_bits_in1,
    output[63:0] mainOff_sub1_req_bits_in2,
    output[9:0] mainOff_sub1_req_tag,
    output mainOff_sub1_rep_ready,
    input  mainOff_sub1_rep_valid,
    input [63:0] mainOff_sub1_rep_bits_out,
    input [9:0] mainOff_sub1_rep_tag,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] T0;
  wire[9:0] T1;
  wire T2;
  wire T3;
  wire[1:0] T4;
  wire rThreadEncoder_io_chosen;
  wire T5;
  reg[0:0] subStateTh_0;
  wire T6;
  wire T7;
  wire T8;
  wire vThreadEncoder_io_chosen;
  wire T9;
  wire AllOffloadsValid_0;
  wire T10;
  wire T11;
  wire T12;
  reg[0:0] sqrtPortHadValidRequest_0;
  wire T13;
  wire T14;
  wire T15;
  wire sqrtPort_req_valid;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  reg[7:0] State_0;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[7:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire[7:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire[7:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire sThreadEncoder_io_chosen;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  reg[7:0] EmitReturnState_0;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] sqrt_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] sqrtPort_rep_tag;
  wire sqrtPort_rep_ready;
  wire[9:0] sqrtPort_req_tag;
  wire[9:0] T104;
  wire sqrtPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  reg[0:0] mul3PortHadValidRequest_0;
  wire T121;
  wire T122;
  wire T123;
  wire mul3Port_req_valid;
  wire T124;
  wire T125;
  wire T126;
  wire[7:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] mul3_valid_received_0;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire[9:0] T136;
  wire[9:0] mul3Port_rep_tag;
  wire mul3Port_rep_ready;
  wire[9:0] mul3Port_req_tag;
  wire[9:0] T137;
  wire mul3Port_rep_valid;
  wire T138;
  wire T139;
  wire[4:0] T140;
  wire T141;
  wire T142;
  wire[4:0] T143;
  wire T144;
  wire T145;
  wire[4:0] T146;
  wire T147;
  wire T148;
  wire T149;
  wire[9:0] T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] mul2PortHadValidRequest_0;
  wire T154;
  wire T155;
  wire T156;
  wire mul2Port_req_valid;
  wire T157;
  wire T158;
  wire T159;
  wire[7:0] T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  reg[0:0] mul2_valid_received_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire[9:0] T169;
  wire[9:0] mul2Port_rep_tag;
  wire mul2Port_rep_ready;
  wire[9:0] mul2Port_req_tag;
  wire[9:0] T170;
  wire mul2Port_rep_valid;
  wire T171;
  wire T172;
  wire[4:0] T173;
  wire T174;
  wire T175;
  wire[4:0] T176;
  wire T177;
  wire T178;
  wire[4:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire[9:0] T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] mul1PortHadValidRequest_0;
  wire T187;
  wire T188;
  wire T189;
  wire mul1Port_req_valid;
  wire T190;
  wire T191;
  wire T192;
  wire[7:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] mul1_valid_received_0;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[9:0] T202;
  wire[9:0] mul1Port_rep_tag;
  wire mul1Port_rep_ready;
  wire[9:0] mul1Port_req_tag;
  wire[9:0] T203;
  wire mul1Port_rep_valid;
  wire T204;
  wire T205;
  wire[4:0] T206;
  wire T207;
  wire T208;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire[4:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[9:0] T216;
  wire T217;
  wire T218;
  wire T219;
  reg[0:0] add2PortHadValidRequest_0;
  wire T220;
  wire T221;
  wire T222;
  wire add2Port_req_valid;
  wire T223;
  wire T224;
  wire T225;
  wire[7:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  reg[0:0] add2_valid_received_0;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[9:0] T235;
  wire[9:0] add2Port_rep_tag;
  wire add2Port_rep_ready;
  wire[9:0] add2Port_req_tag;
  wire[9:0] T236;
  wire add2Port_rep_valid;
  wire T237;
  wire T238;
  wire[4:0] T239;
  wire T240;
  wire T241;
  wire[4:0] T242;
  wire T243;
  wire T244;
  wire[4:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[9:0] T249;
  wire T250;
  wire T251;
  wire T252;
  reg[0:0] add1PortHadValidRequest_0;
  wire T253;
  wire T254;
  wire T255;
  wire add1Port_req_valid;
  wire T256;
  wire T257;
  wire T258;
  wire[7:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg[0:0] add1_valid_received_0;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[9:0] T268;
  wire[9:0] add1Port_rep_tag;
  wire add1Port_rep_ready;
  wire[9:0] add1Port_req_tag;
  wire[9:0] T269;
  wire add1Port_rep_valid;
  wire T270;
  wire T271;
  wire[4:0] T272;
  wire T273;
  wire T274;
  wire[4:0] T275;
  wire T276;
  wire T277;
  wire[4:0] T278;
  wire T279;
  wire T280;
  wire T281;
  wire[9:0] T282;
  wire T283;
  wire T284;
  wire T285;
  reg[0:0] sub3PortHadValidRequest_0;
  wire T286;
  wire T287;
  wire T288;
  wire sub3Port_req_valid;
  wire T289;
  wire T290;
  wire T291;
  wire[7:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  reg[0:0] sub3_valid_received_0;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire[9:0] T301;
  wire[9:0] sub3Port_rep_tag;
  wire sub3Port_rep_ready;
  wire[9:0] sub3Port_req_tag;
  wire[9:0] T302;
  wire sub3Port_rep_valid;
  wire T303;
  wire T304;
  wire[4:0] T305;
  wire T306;
  wire T307;
  wire[4:0] T308;
  wire T309;
  wire T310;
  wire[4:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[9:0] T315;
  wire T316;
  wire T317;
  wire T318;
  reg[0:0] sub2PortHadValidRequest_0;
  wire T319;
  wire T320;
  wire T321;
  wire sub2Port_req_valid;
  wire T322;
  wire T323;
  wire T324;
  wire[7:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  reg[0:0] sub2_valid_received_0;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire[9:0] T334;
  wire[9:0] sub2Port_rep_tag;
  wire sub2Port_rep_ready;
  wire[9:0] sub2Port_req_tag;
  wire[9:0] T335;
  wire sub2Port_rep_valid;
  wire T336;
  wire T337;
  wire[4:0] T338;
  wire T339;
  wire T340;
  wire[4:0] T341;
  wire T342;
  wire T343;
  wire[4:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[9:0] T348;
  wire T349;
  wire T350;
  reg[0:0] sub1PortHadValidRequest_0;
  wire T351;
  wire T352;
  wire T353;
  wire sub1Port_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire[7:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg[0:0] sub1_valid_received_0;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire[9:0] T366;
  wire[9:0] sub1Port_rep_tag;
  wire sub1Port_rep_ready;
  wire[9:0] sub1Port_req_tag;
  wire[9:0] T367;
  wire sub1Port_rep_valid;
  wire T368;
  wire T369;
  wire[4:0] T370;
  wire T371;
  wire T372;
  wire[4:0] T373;
  wire T374;
  wire T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire[9:0] T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire AllOffloadsReady;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  reg[0:0] sqrtPortHadReadyRequest;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg[0:0] sqrt_ready_received;
  wire T397;
  wire T398;
  wire sqrtPort_req_ready;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg[0:0] mul3PortHadReadyRequest;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg[0:0] mul3_ready_received;
  wire T409;
  wire T410;
  wire mul3Port_req_ready;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg[0:0] mul2PortHadReadyRequest;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg[0:0] mul2_ready_received;
  wire T421;
  wire T422;
  wire mul2Port_req_ready;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  reg[0:0] mul1PortHadReadyRequest;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg[0:0] mul1_ready_received;
  wire T433;
  wire T434;
  wire mul1Port_req_ready;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  reg[0:0] add2PortHadReadyRequest;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg[0:0] add2_ready_received;
  wire T445;
  wire T446;
  wire add2Port_req_ready;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  reg[0:0] add1PortHadReadyRequest;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg[0:0] add1_ready_received;
  wire T457;
  wire T458;
  wire add1Port_req_ready;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  reg[0:0] sub3PortHadReadyRequest;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  reg[0:0] sub3_ready_received;
  wire T469;
  wire T470;
  wire sub3Port_req_ready;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  reg[0:0] sub2PortHadReadyRequest;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  reg[0:0] sub2_ready_received;
  wire T481;
  wire T482;
  wire sub2Port_req_ready;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg[0:0] sub1PortHadReadyRequest;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  reg[0:0] sub1_ready_received;
  wire T492;
  wire T493;
  wire sub1Port_req_ready;
  wire T494;
  reg[9:0] inputTag_0;
  wire[9:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;

  assign io_out_tag = T0;
  assign T0 = inputTag_0 & T1;
  assign T1 = {4'ha/* 10*/{T2}};
  assign T2 = T3;
  assign T3 = T4[1'h0/* 0*/:1'h0/* 0*/];
  assign T4 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T5 = subStateTh_0 == 1'h0/* 0*/;
  assign T6 = T382 ? 1'h1/* 1*/ : T7;
  assign T7 = T8 ? 1'h0/* 0*/ : subStateTh_0;
  assign T8 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T9 = T381 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T10;
  assign T10 = T118 && T11;
  assign T11 = T114 || T12;
  assign T12 = ! sqrtPortHadValidRequest_0;
  assign T13 = T111 && T14;
  assign T14 = sqrtPortHadValidRequest_0 || T15;
  assign T15 = T109 && sqrtPort_req_valid;
  assign sqrtPort_req_valid = T16;
  assign T16 = T96 && T17;
  assign T17 = T95 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T2}};
  assign T22 = T33 || T23;
  assign T23 = T27 && T24;
  assign T24 = T25;
  assign T25 = T26[1'h0/* 0*/:1'h0/* 0*/];
  assign T26 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T27 = T32 && T28;
  assign T28 = T30 == T29;
  assign T29 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T30 = State_0 & T31;
  assign T31 = {4'h8/* 8*/{T24}};
  assign T32 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T33 = T39 || T34;
  assign T34 = T35 && T24;
  assign T35 = T38 && T36;
  assign T36 = T30 == T37;
  assign T37 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T38 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T39 = T45 || T40;
  assign T40 = T41 && T24;
  assign T41 = T44 && T42;
  assign T42 = T30 == T43;
  assign T43 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T44 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T45 = T51 || T46;
  assign T46 = T47 && T24;
  assign T47 = T50 && T48;
  assign T48 = T30 == T49;
  assign T49 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T50 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T51 = T57 || T52;
  assign T52 = T53 && T24;
  assign T53 = T56 && T54;
  assign T54 = T30 == T55;
  assign T55 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T56 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T57 = T63 || T58;
  assign T58 = T59 && T24;
  assign T59 = T62 && T60;
  assign T60 = T30 == T61;
  assign T61 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T62 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T63 = T69 || T64;
  assign T64 = T65 && T2;
  assign T65 = T66 && io_out_ready;
  assign T66 = T68 && T67;
  assign T67 = T20 == 8'hff/* 255*/;
  assign T68 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T69 = T76 && T70;
  assign T70 = T71;
  assign T71 = T72[1'h0/* 0*/:1'h0/* 0*/];
  assign T72 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T73 = T75 && T74;
  assign T74 = State_0 == 8'h0/* 0*/;
  assign T75 = subStateTh_0 == 1'h0/* 0*/;
  assign T76 = T77 && io_in_valid;
  assign T77 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = T23 ? 8'hff/* 255*/ : T79;
  assign T79 = T34 ? T94 : T80;
  assign T80 = T40 ? T93 : T81;
  assign T81 = T46 ? T92 : T82;
  assign T82 = T52 ? T91 : T83;
  assign T83 = T58 ? T90 : T84;
  assign T84 = T64 ? T87 : T85;
  assign T85 = T69 ? T86 : State_0;
  assign T86 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T87 = EmitReturnState_0 & T88;
  assign T88 = {4'h8/* 8*/{T2}};
  assign T89 = T23 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T90 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T91 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T92 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T93 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T94 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = sqrt_valid_received_0 & T2;
  assign T99 = T105 && T100;
  assign T100 = sqrt_valid_received_0 || T101;
  assign T101 = sqrtPort_rep_valid && T102;
  assign T102 = sqrtPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sqrtPort_rep_tag = mainOff_sqrt_rep_tag;
  assign mainOff_sqrt_rep_ready = sqrtPort_rep_ready;
  assign sqrtPort_rep_ready = 1'h1/* 1*/;
  assign mainOff_sqrt_req_tag = sqrtPort_req_tag;
  assign sqrtPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sqrtPort_rep_valid = mainOff_sqrt_rep_valid;
  assign mainOff_sqrt_req_valid = sqrtPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || sqrt_valid_received_0;
  assign T115 = sqrtPort_rep_valid && T116;
  assign T116 = sqrtPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T151 && T119;
  assign T119 = T147 || T120;
  assign T120 = ! mul3PortHadValidRequest_0;
  assign T121 = T144 && T122;
  assign T122 = mul3PortHadValidRequest_0 || T123;
  assign T123 = T142 && mul3Port_req_valid;
  assign mul3Port_req_valid = T124;
  assign T124 = T129 && T125;
  assign T125 = T128 && T126;
  assign T126 = T20 == T127;
  assign T127 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T128 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T129 = T141 && T130;
  assign T130 = ! T131;
  assign T131 = mul3_valid_received_0 & T2;
  assign T132 = T138 && T133;
  assign T133 = mul3_valid_received_0 || T134;
  assign T134 = mul3Port_rep_valid && T135;
  assign T135 = mul3Port_rep_tag == T136;
  assign T136 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul3Port_rep_tag = mainOff_mul3_rep_tag;
  assign mainOff_mul3_rep_ready = mul3Port_rep_ready;
  assign mul3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul3_req_tag = mul3Port_req_tag;
  assign mul3Port_req_tag = T137;
  assign T137 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul3Port_rep_valid = mainOff_mul3_rep_valid;
  assign mainOff_mul3_req_valid = mul3Port_req_valid;
  assign T138 = ! T139;
  assign T139 = T140 == 5'h0/* 0*/;
  assign T140 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T141 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T142 = 5'h0/* 0*/ == T143;
  assign T143 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T144 = ! T145;
  assign T145 = T146 == 5'h0/* 0*/;
  assign T146 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T147 = T148 || mul3_valid_received_0;
  assign T148 = mul3Port_rep_valid && T149;
  assign T149 = mul3Port_rep_tag == T150;
  assign T150 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T151 = T184 && T152;
  assign T152 = T180 || T153;
  assign T153 = ! mul2PortHadValidRequest_0;
  assign T154 = T177 && T155;
  assign T155 = mul2PortHadValidRequest_0 || T156;
  assign T156 = T175 && mul2Port_req_valid;
  assign mul2Port_req_valid = T157;
  assign T157 = T162 && T158;
  assign T158 = T161 && T159;
  assign T159 = T20 == T160;
  assign T160 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T161 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T162 = T174 && T163;
  assign T163 = ! T164;
  assign T164 = mul2_valid_received_0 & T2;
  assign T165 = T171 && T166;
  assign T166 = mul2_valid_received_0 || T167;
  assign T167 = mul2Port_rep_valid && T168;
  assign T168 = mul2Port_rep_tag == T169;
  assign T169 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul2Port_rep_tag = mainOff_mul2_rep_tag;
  assign mainOff_mul2_rep_ready = mul2Port_rep_ready;
  assign mul2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul2_req_tag = mul2Port_req_tag;
  assign mul2Port_req_tag = T170;
  assign T170 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul2Port_rep_valid = mainOff_mul2_rep_valid;
  assign mainOff_mul2_req_valid = mul2Port_req_valid;
  assign T171 = ! T172;
  assign T172 = T173 == 5'h0/* 0*/;
  assign T173 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T174 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T175 = 5'h0/* 0*/ == T176;
  assign T176 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T177 = ! T178;
  assign T178 = T179 == 5'h0/* 0*/;
  assign T179 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T180 = T181 || mul2_valid_received_0;
  assign T181 = mul2Port_rep_valid && T182;
  assign T182 = mul2Port_rep_tag == T183;
  assign T183 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T184 = T217 && T185;
  assign T185 = T213 || T186;
  assign T186 = ! mul1PortHadValidRequest_0;
  assign T187 = T210 && T188;
  assign T188 = mul1PortHadValidRequest_0 || T189;
  assign T189 = T208 && mul1Port_req_valid;
  assign mul1Port_req_valid = T190;
  assign T190 = T195 && T191;
  assign T191 = T194 && T192;
  assign T192 = T20 == T193;
  assign T193 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T194 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T195 = T207 && T196;
  assign T196 = ! T197;
  assign T197 = mul1_valid_received_0 & T2;
  assign T198 = T204 && T199;
  assign T199 = mul1_valid_received_0 || T200;
  assign T200 = mul1Port_rep_valid && T201;
  assign T201 = mul1Port_rep_tag == T202;
  assign T202 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign mul1Port_rep_tag = mainOff_mul1_rep_tag;
  assign mainOff_mul1_rep_ready = mul1Port_rep_ready;
  assign mul1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_mul1_req_tag = mul1Port_req_tag;
  assign mul1Port_req_tag = T203;
  assign T203 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign mul1Port_rep_valid = mainOff_mul1_rep_valid;
  assign mainOff_mul1_req_valid = mul1Port_req_valid;
  assign T204 = ! T205;
  assign T205 = T206 == 5'h0/* 0*/;
  assign T206 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T207 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T208 = 5'h0/* 0*/ == T209;
  assign T209 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T210 = ! T211;
  assign T211 = T212 == 5'h0/* 0*/;
  assign T212 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T213 = T214 || mul1_valid_received_0;
  assign T214 = mul1Port_rep_valid && T215;
  assign T215 = mul1Port_rep_tag == T216;
  assign T216 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T217 = T250 && T218;
  assign T218 = T246 || T219;
  assign T219 = ! add2PortHadValidRequest_0;
  assign T220 = T243 && T221;
  assign T221 = add2PortHadValidRequest_0 || T222;
  assign T222 = T241 && add2Port_req_valid;
  assign add2Port_req_valid = T223;
  assign T223 = T228 && T224;
  assign T224 = T227 && T225;
  assign T225 = T20 == T226;
  assign T226 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T228 = T240 && T229;
  assign T229 = ! T230;
  assign T230 = add2_valid_received_0 & T2;
  assign T231 = T237 && T232;
  assign T232 = add2_valid_received_0 || T233;
  assign T233 = add2Port_rep_valid && T234;
  assign T234 = add2Port_rep_tag == T235;
  assign T235 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add2Port_rep_tag = mainOff_add2_rep_tag;
  assign mainOff_add2_rep_ready = add2Port_rep_ready;
  assign add2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add2_req_tag = add2Port_req_tag;
  assign add2Port_req_tag = T236;
  assign T236 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add2Port_rep_valid = mainOff_add2_rep_valid;
  assign mainOff_add2_req_valid = add2Port_req_valid;
  assign T237 = ! T238;
  assign T238 = T239 == 5'h0/* 0*/;
  assign T239 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T240 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T241 = 5'h0/* 0*/ == T242;
  assign T242 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T243 = ! T244;
  assign T244 = T245 == 5'h0/* 0*/;
  assign T245 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T246 = T247 || add2_valid_received_0;
  assign T247 = add2Port_rep_valid && T248;
  assign T248 = add2Port_rep_tag == T249;
  assign T249 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T250 = T283 && T251;
  assign T251 = T279 || T252;
  assign T252 = ! add1PortHadValidRequest_0;
  assign T253 = T276 && T254;
  assign T254 = add1PortHadValidRequest_0 || T255;
  assign T255 = T274 && add1Port_req_valid;
  assign add1Port_req_valid = T256;
  assign T256 = T261 && T257;
  assign T257 = T260 && T258;
  assign T258 = T20 == T259;
  assign T259 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T260 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T261 = T273 && T262;
  assign T262 = ! T263;
  assign T263 = add1_valid_received_0 & T2;
  assign T264 = T270 && T265;
  assign T265 = add1_valid_received_0 || T266;
  assign T266 = add1Port_rep_valid && T267;
  assign T267 = add1Port_rep_tag == T268;
  assign T268 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign add1Port_rep_tag = mainOff_add1_rep_tag;
  assign mainOff_add1_rep_ready = add1Port_rep_ready;
  assign add1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_add1_req_tag = add1Port_req_tag;
  assign add1Port_req_tag = T269;
  assign T269 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign add1Port_rep_valid = mainOff_add1_rep_valid;
  assign mainOff_add1_req_valid = add1Port_req_valid;
  assign T270 = ! T271;
  assign T271 = T272 == 5'h0/* 0*/;
  assign T272 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T273 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T274 = 5'h0/* 0*/ == T275;
  assign T275 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T276 = ! T277;
  assign T277 = T278 == 5'h0/* 0*/;
  assign T278 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T279 = T280 || add1_valid_received_0;
  assign T280 = add1Port_rep_valid && T281;
  assign T281 = add1Port_rep_tag == T282;
  assign T282 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T283 = T316 && T284;
  assign T284 = T312 || T285;
  assign T285 = ! sub3PortHadValidRequest_0;
  assign T286 = T309 && T287;
  assign T287 = sub3PortHadValidRequest_0 || T288;
  assign T288 = T307 && sub3Port_req_valid;
  assign sub3Port_req_valid = T289;
  assign T289 = T294 && T290;
  assign T290 = T293 && T291;
  assign T291 = T20 == T292;
  assign T292 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T293 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T294 = T306 && T295;
  assign T295 = ! T296;
  assign T296 = sub3_valid_received_0 & T2;
  assign T297 = T303 && T298;
  assign T298 = sub3_valid_received_0 || T299;
  assign T299 = sub3Port_rep_valid && T300;
  assign T300 = sub3Port_rep_tag == T301;
  assign T301 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub3Port_rep_tag = mainOff_sub3_rep_tag;
  assign mainOff_sub3_rep_ready = sub3Port_rep_ready;
  assign sub3Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub3_req_tag = sub3Port_req_tag;
  assign sub3Port_req_tag = T302;
  assign T302 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub3Port_rep_valid = mainOff_sub3_rep_valid;
  assign mainOff_sub3_req_valid = sub3Port_req_valid;
  assign T303 = ! T304;
  assign T304 = T305 == 5'h0/* 0*/;
  assign T305 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T306 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T307 = 5'h0/* 0*/ == T308;
  assign T308 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T309 = ! T310;
  assign T310 = T311 == 5'h0/* 0*/;
  assign T311 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T312 = T313 || sub3_valid_received_0;
  assign T313 = sub3Port_rep_valid && T314;
  assign T314 = sub3Port_rep_tag == T315;
  assign T315 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T316 = T349 && T317;
  assign T317 = T345 || T318;
  assign T318 = ! sub2PortHadValidRequest_0;
  assign T319 = T342 && T320;
  assign T320 = sub2PortHadValidRequest_0 || T321;
  assign T321 = T340 && sub2Port_req_valid;
  assign sub2Port_req_valid = T322;
  assign T322 = T327 && T323;
  assign T323 = T326 && T324;
  assign T324 = T20 == T325;
  assign T325 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T326 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T327 = T339 && T328;
  assign T328 = ! T329;
  assign T329 = sub2_valid_received_0 & T2;
  assign T330 = T336 && T331;
  assign T331 = sub2_valid_received_0 || T332;
  assign T332 = sub2Port_rep_valid && T333;
  assign T333 = sub2Port_rep_tag == T334;
  assign T334 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub2Port_rep_tag = mainOff_sub2_rep_tag;
  assign mainOff_sub2_rep_ready = sub2Port_rep_ready;
  assign sub2Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub2_req_tag = sub2Port_req_tag;
  assign sub2Port_req_tag = T335;
  assign T335 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub2Port_rep_valid = mainOff_sub2_rep_valid;
  assign mainOff_sub2_req_valid = sub2Port_req_valid;
  assign T336 = ! T337;
  assign T337 = T338 == 5'h0/* 0*/;
  assign T338 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T339 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T340 = 5'h0/* 0*/ == T341;
  assign T341 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T342 = ! T343;
  assign T343 = T344 == 5'h0/* 0*/;
  assign T344 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T345 = T346 || sub2_valid_received_0;
  assign T346 = sub2Port_rep_valid && T347;
  assign T347 = sub2Port_rep_tag == T348;
  assign T348 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T349 = T377 || T350;
  assign T350 = ! sub1PortHadValidRequest_0;
  assign T351 = T374 && T352;
  assign T352 = sub1PortHadValidRequest_0 || T353;
  assign T353 = T372 && sub1Port_req_valid;
  assign sub1Port_req_valid = T354;
  assign T354 = T359 && T355;
  assign T355 = T358 && T356;
  assign T356 = T20 == T357;
  assign T357 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T358 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T359 = T371 && T360;
  assign T360 = ! T361;
  assign T361 = sub1_valid_received_0 & T2;
  assign T362 = T368 && T363;
  assign T363 = sub1_valid_received_0 || T364;
  assign T364 = sub1Port_rep_valid && T365;
  assign T365 = sub1Port_rep_tag == T366;
  assign T366 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign sub1Port_rep_tag = mainOff_sub1_rep_tag;
  assign mainOff_sub1_rep_ready = sub1Port_rep_ready;
  assign sub1Port_rep_ready = 1'h1/* 1*/;
  assign mainOff_sub1_req_tag = sub1Port_req_tag;
  assign sub1Port_req_tag = T367;
  assign T367 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign sub1Port_rep_valid = mainOff_sub1_rep_valid;
  assign mainOff_sub1_req_valid = sub1Port_req_valid;
  assign T368 = ! T369;
  assign T369 = T370 == 5'h0/* 0*/;
  assign T370 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T371 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T372 = 5'h0/* 0*/ == T373;
  assign T373 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T374 = ! T375;
  assign T375 = T376 == 5'h0/* 0*/;
  assign T376 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T377 = T378 || sub1_valid_received_0;
  assign T378 = sub1Port_rep_valid && T379;
  assign T379 = sub1Port_rep_tag == T380;
  assign T380 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T381 = subStateTh_0 == 1'h1/* 1*/;
  assign T382 = T384 && T383;
  assign T383 = State_0 != 8'hff/* 255*/;
  assign T384 = T386 && T385;
  assign T385 = State_0 != 8'h0/* 0*/;
  assign T386 = AllOffloadsReady && T387;
  assign T387 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T388;
  assign T388 = T400 && T389;
  assign T389 = T396 || T390;
  assign T390 = T392 && T391;
  assign T391 = ! sqrtPort_req_valid;
  assign T392 = ! sqrtPortHadReadyRequest;
  assign T393 = T395 && T394;
  assign T394 = sqrtPortHadReadyRequest || sqrtPort_req_valid;
  assign T395 = ! AllOffloadsReady;
  assign T396 = sqrtPort_req_ready || sqrt_ready_received;
  assign T397 = T399 && T398;
  assign T398 = sqrt_ready_received || sqrtPort_req_ready;
  assign sqrtPort_req_ready = mainOff_sqrt_req_ready;
  assign T399 = ! AllOffloadsReady;
  assign T400 = T412 && T401;
  assign T401 = T408 || T402;
  assign T402 = T404 && T403;
  assign T403 = ! mul3Port_req_valid;
  assign T404 = ! mul3PortHadReadyRequest;
  assign T405 = T407 && T406;
  assign T406 = mul3PortHadReadyRequest || mul3Port_req_valid;
  assign T407 = ! AllOffloadsReady;
  assign T408 = mul3Port_req_ready || mul3_ready_received;
  assign T409 = T411 && T410;
  assign T410 = mul3_ready_received || mul3Port_req_ready;
  assign mul3Port_req_ready = mainOff_mul3_req_ready;
  assign T411 = ! AllOffloadsReady;
  assign T412 = T424 && T413;
  assign T413 = T420 || T414;
  assign T414 = T416 && T415;
  assign T415 = ! mul2Port_req_valid;
  assign T416 = ! mul2PortHadReadyRequest;
  assign T417 = T419 && T418;
  assign T418 = mul2PortHadReadyRequest || mul2Port_req_valid;
  assign T419 = ! AllOffloadsReady;
  assign T420 = mul2Port_req_ready || mul2_ready_received;
  assign T421 = T423 && T422;
  assign T422 = mul2_ready_received || mul2Port_req_ready;
  assign mul2Port_req_ready = mainOff_mul2_req_ready;
  assign T423 = ! AllOffloadsReady;
  assign T424 = T436 && T425;
  assign T425 = T432 || T426;
  assign T426 = T428 && T427;
  assign T427 = ! mul1Port_req_valid;
  assign T428 = ! mul1PortHadReadyRequest;
  assign T429 = T431 && T430;
  assign T430 = mul1PortHadReadyRequest || mul1Port_req_valid;
  assign T431 = ! AllOffloadsReady;
  assign T432 = mul1Port_req_ready || mul1_ready_received;
  assign T433 = T435 && T434;
  assign T434 = mul1_ready_received || mul1Port_req_ready;
  assign mul1Port_req_ready = mainOff_mul1_req_ready;
  assign T435 = ! AllOffloadsReady;
  assign T436 = T448 && T437;
  assign T437 = T444 || T438;
  assign T438 = T440 && T439;
  assign T439 = ! add2Port_req_valid;
  assign T440 = ! add2PortHadReadyRequest;
  assign T441 = T443 && T442;
  assign T442 = add2PortHadReadyRequest || add2Port_req_valid;
  assign T443 = ! AllOffloadsReady;
  assign T444 = add2Port_req_ready || add2_ready_received;
  assign T445 = T447 && T446;
  assign T446 = add2_ready_received || add2Port_req_ready;
  assign add2Port_req_ready = mainOff_add2_req_ready;
  assign T447 = ! AllOffloadsReady;
  assign T448 = T460 && T449;
  assign T449 = T456 || T450;
  assign T450 = T452 && T451;
  assign T451 = ! add1Port_req_valid;
  assign T452 = ! add1PortHadReadyRequest;
  assign T453 = T455 && T454;
  assign T454 = add1PortHadReadyRequest || add1Port_req_valid;
  assign T455 = ! AllOffloadsReady;
  assign T456 = add1Port_req_ready || add1_ready_received;
  assign T457 = T459 && T458;
  assign T458 = add1_ready_received || add1Port_req_ready;
  assign add1Port_req_ready = mainOff_add1_req_ready;
  assign T459 = ! AllOffloadsReady;
  assign T460 = T472 && T461;
  assign T461 = T468 || T462;
  assign T462 = T464 && T463;
  assign T463 = ! sub3Port_req_valid;
  assign T464 = ! sub3PortHadReadyRequest;
  assign T465 = T467 && T466;
  assign T466 = sub3PortHadReadyRequest || sub3Port_req_valid;
  assign T467 = ! AllOffloadsReady;
  assign T468 = sub3Port_req_ready || sub3_ready_received;
  assign T469 = T471 && T470;
  assign T470 = sub3_ready_received || sub3Port_req_ready;
  assign sub3Port_req_ready = mainOff_sub3_req_ready;
  assign T471 = ! AllOffloadsReady;
  assign T472 = T484 && T473;
  assign T473 = T480 || T474;
  assign T474 = T476 && T475;
  assign T475 = ! sub2Port_req_valid;
  assign T476 = ! sub2PortHadReadyRequest;
  assign T477 = T479 && T478;
  assign T478 = sub2PortHadReadyRequest || sub2Port_req_valid;
  assign T479 = ! AllOffloadsReady;
  assign T480 = sub2Port_req_ready || sub2_ready_received;
  assign T481 = T483 && T482;
  assign T482 = sub2_ready_received || sub2Port_req_ready;
  assign sub2Port_req_ready = mainOff_sub2_req_ready;
  assign T483 = ! AllOffloadsReady;
  assign T484 = T491 || T485;
  assign T485 = T487 && T486;
  assign T486 = ! sub1Port_req_valid;
  assign T487 = ! sub1PortHadReadyRequest;
  assign T488 = T490 && T489;
  assign T489 = sub1PortHadReadyRequest || sub1Port_req_valid;
  assign T490 = ! AllOffloadsReady;
  assign T491 = sub1Port_req_ready || sub1_ready_received;
  assign T492 = T494 && T493;
  assign T493 = sub1_ready_received || sub1Port_req_ready;
  assign sub1Port_req_ready = mainOff_sub1_req_ready;
  assign T494 = ! AllOffloadsReady;
  assign T495 = T69 ? io_in_tag : inputTag_0;
  assign io_out_valid = T496;
  assign T496 = T498 && T497;
  assign T497 = T20 == 8'hff/* 255*/;
  assign T498 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_in_ready = T499;
  assign T499 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  RREncode_60 rThreadEncoder(
       .io_valid_0( T5 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_61 vThreadEncoder(
       .io_valid_0( T9 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_62 sThreadEncoder(
       .io_valid_0( T73 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T6;
    sqrtPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T13;
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T22) begin
      State_0 <= T78;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T23) begin
      EmitReturnState_0 <= T89;
    end
    sqrt_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    mul3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T121;
    mul3_valid_received_0 <= reset ? 1'h0/* 0*/ : T132;
    mul2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T154;
    mul2_valid_received_0 <= reset ? 1'h0/* 0*/ : T165;
    mul1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T187;
    mul1_valid_received_0 <= reset ? 1'h0/* 0*/ : T198;
    add2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T220;
    add2_valid_received_0 <= reset ? 1'h0/* 0*/ : T231;
    add1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T253;
    add1_valid_received_0 <= reset ? 1'h0/* 0*/ : T264;
    sub3PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T286;
    sub3_valid_received_0 <= reset ? 1'h0/* 0*/ : T297;
    sub2PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T319;
    sub2_valid_received_0 <= reset ? 1'h0/* 0*/ : T330;
    sub1PortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T351;
    sub1_valid_received_0 <= reset ? 1'h0/* 0*/ : T362;
    sqrtPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T393;
    sqrt_ready_received <= reset ? 1'h0/* 0*/ : T397;
    mul3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T405;
    mul3_ready_received <= reset ? 1'h0/* 0*/ : T409;
    mul2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T417;
    mul2_ready_received <= reset ? 1'h0/* 0*/ : T421;
    mul1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T429;
    mul1_ready_received <= reset ? 1'h0/* 0*/ : T433;
    add2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T441;
    add2_ready_received <= reset ? 1'h0/* 0*/ : T445;
    add1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T453;
    add1_ready_received <= reset ? 1'h0/* 0*/ : T457;
    sub3PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T465;
    sub3_ready_received <= reset ? 1'h0/* 0*/ : T469;
    sub2PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T477;
    sub2_ready_received <= reset ? 1'h0/* 0*/ : T481;
    sub1PortHadReadyRequest <= reset ? 1'h0/* 0*/ : T488;
    sub1_ready_received <= reset ? 1'h0/* 0*/ : T492;
    if(T69) begin
      inputTag_0 <= T495;
    end
  end
endmodule

module gPipe_90(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_90(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_90 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_117(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub2_req_ready,
    output mainOff_sub2_req_valid,
    output[63:0] mainOff_sub2_req_bits_in1,
    output[63:0] mainOff_sub2_req_bits_in2,
    output[9:0] mainOff_sub2_req_tag,
    output mainOff_sub2_rep_ready,
    input  mainOff_sub2_rep_valid,
    input [63:0] mainOff_sub2_rep_bits_out,
    input [9:0] mainOff_sub2_rep_tag,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire mainComp_mainOff_sub2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub1_rep_ready;
  wire[9:0] mainComp_mainOff_sub1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign mainOff_sub2_rep_ready = mainComp_mainOff_sub2_rep_ready;
  assign mainOff_sub2_req_tag = mainComp_mainOff_sub2_req_tag;
  assign mainOff_sub2_req_valid = mainComp_mainOff_sub2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  distanceFU_9 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y(  ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y(  ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub1_req_ready( offComp_io_in_ready ),
       .mainOff_sub1_req_valid( mainComp_mainOff_sub1_req_valid ),
       .mainOff_sub1_req_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .mainOff_sub1_req_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .mainOff_sub1_req_tag( mainComp_mainOff_sub1_req_tag ),
       .mainOff_sub1_rep_ready( mainComp_mainOff_sub1_rep_ready ),
       .mainOff_sub1_rep_valid( offComp_io_out_valid ),
       .mainOff_sub1_rep_bits_out(  ),
       .mainOff_sub1_rep_tag( offComp_io_out_tag ),
       .mainOff_sub2_req_ready( mainOff_sub2_req_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1(  ),
       .mainOff_sub2_req_bits_in2(  ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( mainOff_sub2_rep_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( mainOff_sub2_rep_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_90 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub1_req_tag ),
       .io_out_ready( mainComp_mainOff_sub1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_91(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_91(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_91 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_118(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sub3_req_ready,
    output mainOff_sub3_req_valid,
    output[63:0] mainOff_sub3_req_bits_in1,
    output[63:0] mainOff_sub3_req_bits_in2,
    output[9:0] mainOff_sub3_req_tag,
    output mainOff_sub3_rep_ready,
    input  mainOff_sub3_rep_valid,
    input [63:0] mainOff_sub3_rep_bits_out,
    input [9:0] mainOff_sub3_rep_tag,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire mainComp_mainOff_sub3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub2_rep_ready;
  wire[9:0] mainComp_mainOff_sub2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign mainOff_sub3_rep_ready = mainComp_mainOff_sub3_rep_ready;
  assign mainOff_sub3_req_tag = mainComp_mainOff_sub3_req_tag;
  assign mainOff_sub3_req_valid = mainComp_mainOff_sub3_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_117 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z(  ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub2_req_ready( offComp_io_in_ready ),
       .mainOff_sub2_req_valid( mainComp_mainOff_sub2_req_valid ),
       .mainOff_sub2_req_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .mainOff_sub2_req_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .mainOff_sub2_req_tag( mainComp_mainOff_sub2_req_tag ),
       .mainOff_sub2_rep_ready( mainComp_mainOff_sub2_rep_ready ),
       .mainOff_sub2_rep_valid( offComp_io_out_valid ),
       .mainOff_sub2_rep_bits_out(  ),
       .mainOff_sub2_rep_tag( offComp_io_out_tag ),
       .mainOff_sub3_req_ready( mainOff_sub3_req_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1(  ),
       .mainOff_sub3_req_bits_in2(  ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( mainOff_sub3_rep_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( mainOff_sub3_rep_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_91 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub2_req_tag ),
       .io_out_ready( mainComp_mainOff_sub2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_92(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_92(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_92 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_119(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul1_req_ready,
    output mainOff_mul1_req_valid,
    output[63:0] mainOff_mul1_req_bits_in1,
    output[63:0] mainOff_mul1_req_bits_in2,
    output[9:0] mainOff_mul1_req_tag,
    output mainOff_mul1_rep_ready,
    input  mainOff_mul1_rep_valid,
    input [63:0] mainOff_mul1_rep_bits_out,
    input [9:0] mainOff_mul1_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sub3_rep_ready;
  wire[9:0] mainComp_mainOff_sub3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sub3_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in1;
  wire[63:0] mainComp_mainOff_sub3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_mul1_rep_ready = mainComp_mainOff_mul1_rep_ready;
  assign mainOff_mul1_req_tag = mainComp_mainOff_mul1_req_tag;
  assign mainOff_mul1_req_valid = mainComp_mainOff_mul1_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_118 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sub3_req_ready( offComp_io_in_ready ),
       .mainOff_sub3_req_valid( mainComp_mainOff_sub3_req_valid ),
       .mainOff_sub3_req_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .mainOff_sub3_req_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .mainOff_sub3_req_tag( mainComp_mainOff_sub3_req_tag ),
       .mainOff_sub3_rep_ready( mainComp_mainOff_sub3_rep_ready ),
       .mainOff_sub3_rep_valid( offComp_io_out_valid ),
       .mainOff_sub3_rep_bits_out(  ),
       .mainOff_sub3_rep_tag( offComp_io_out_tag ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( mainOff_mul1_req_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1(  ),
       .mainOff_mul1_req_bits_in2(  ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( mainOff_mul1_rep_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( mainOff_mul1_rep_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_92 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sub3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sub3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sub3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sub3_req_tag ),
       .io_out_ready( mainComp_mainOff_sub3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_93(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_93(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_93 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_120(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul2_req_ready,
    output mainOff_mul2_req_valid,
    output[63:0] mainOff_mul2_req_bits_in1,
    output[63:0] mainOff_mul2_req_bits_in2,
    output[9:0] mainOff_mul2_req_tag,
    output mainOff_mul2_rep_ready,
    input  mainOff_mul2_rep_valid,
    input [63:0] mainOff_mul2_rep_bits_out,
    input [9:0] mainOff_mul2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire mainComp_mainOff_mul2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul1_rep_ready;
  wire[9:0] mainComp_mainOff_mul1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul1_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_mul2_rep_ready = mainComp_mainOff_mul2_rep_ready;
  assign mainOff_mul2_req_tag = mainComp_mainOff_mul2_req_tag;
  assign mainOff_mul2_req_valid = mainComp_mainOff_mul2_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_119 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul1_req_ready( offComp_io_in_ready ),
       .mainOff_mul1_req_valid( mainComp_mainOff_mul1_req_valid ),
       .mainOff_mul1_req_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .mainOff_mul1_req_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .mainOff_mul1_req_tag( mainComp_mainOff_mul1_req_tag ),
       .mainOff_mul1_rep_ready( mainComp_mainOff_mul1_rep_ready ),
       .mainOff_mul1_rep_valid( offComp_io_out_valid ),
       .mainOff_mul1_rep_bits_out(  ),
       .mainOff_mul1_rep_tag( offComp_io_out_tag ),
       .mainOff_mul2_req_ready( mainOff_mul2_req_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1(  ),
       .mainOff_mul2_req_bits_in2(  ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( mainOff_mul2_rep_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( mainOff_mul2_rep_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_93 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul1_req_tag ),
       .io_out_ready( mainComp_mainOff_mul1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_94(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_94(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_94 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_121(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_mul3_req_ready,
    output mainOff_mul3_req_valid,
    output[63:0] mainOff_mul3_req_bits_in1,
    output[63:0] mainOff_mul3_req_bits_in2,
    output[9:0] mainOff_mul3_req_tag,
    output mainOff_mul3_rep_ready,
    input  mainOff_mul3_rep_valid,
    input [63:0] mainOff_mul3_rep_bits_out,
    input [9:0] mainOff_mul3_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire mainComp_mainOff_mul3_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul2_rep_ready;
  wire[9:0] mainComp_mainOff_mul2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul2_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_mul3_rep_ready = mainComp_mainOff_mul3_rep_ready;
  assign mainOff_mul3_req_tag = mainComp_mainOff_mul3_req_tag;
  assign mainOff_mul3_req_valid = mainComp_mainOff_mul3_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_120 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul2_req_ready( offComp_io_in_ready ),
       .mainOff_mul2_req_valid( mainComp_mainOff_mul2_req_valid ),
       .mainOff_mul2_req_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .mainOff_mul2_req_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .mainOff_mul2_req_tag( mainComp_mainOff_mul2_req_tag ),
       .mainOff_mul2_rep_ready( mainComp_mainOff_mul2_rep_ready ),
       .mainOff_mul2_rep_valid( offComp_io_out_valid ),
       .mainOff_mul2_rep_bits_out(  ),
       .mainOff_mul2_rep_tag( offComp_io_out_tag ),
       .mainOff_mul3_req_ready( mainOff_mul3_req_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1(  ),
       .mainOff_mul3_req_bits_in2(  ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( mainOff_mul3_rep_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( mainOff_mul3_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_94 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul2_req_tag ),
       .io_out_ready( mainComp_mainOff_mul2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_95(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_95(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_95 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_93_ACMP_dmul_3_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_122(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add1_req_ready,
    output mainOff_add1_req_valid,
    output[63:0] mainOff_add1_req_bits_in1,
    output[63:0] mainOff_add1_req_bits_in2,
    output[9:0] mainOff_add1_req_tag,
    output mainOff_add1_rep_ready,
    input  mainOff_add1_rep_valid,
    input [63:0] mainOff_add1_rep_bits_out,
    input [9:0] mainOff_add1_rep_tag,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_mul3_rep_ready;
  wire[9:0] mainComp_mainOff_mul3_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_mul3_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in1;
  wire[63:0] mainComp_mainOff_mul3_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign mainOff_add1_rep_ready = mainComp_mainOff_add1_rep_ready;
  assign mainOff_add1_req_tag = mainComp_mainOff_add1_req_tag;
  assign mainOff_add1_req_valid = mainComp_mainOff_add1_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_121 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( mainOff_add1_req_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1(  ),
       .mainOff_add1_req_bits_in2(  ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( mainOff_add1_rep_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( mainOff_add1_rep_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_mul3_req_ready( offComp_io_in_ready ),
       .mainOff_mul3_req_valid( mainComp_mainOff_mul3_req_valid ),
       .mainOff_mul3_req_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .mainOff_mul3_req_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .mainOff_mul3_req_tag( mainComp_mainOff_mul3_req_tag ),
       .mainOff_mul3_rep_ready( mainComp_mainOff_mul3_rep_ready ),
       .mainOff_mul3_rep_valid( offComp_io_out_valid ),
       .mainOff_mul3_rep_bits_out(  ),
       .mainOff_mul3_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_95 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_mul3_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_mul3_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_mul3_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_mul3_req_tag ),
       .io_out_ready( mainComp_mainOff_mul3_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_96(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_96(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_96 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_123(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add2_req_ready,
    output mainOff_add2_req_valid,
    output[63:0] mainOff_add2_req_bits_in1,
    output[63:0] mainOff_add2_req_bits_in2,
    output[9:0] mainOff_add2_req_tag,
    output mainOff_add2_rep_ready,
    input  mainOff_add2_rep_valid,
    input [63:0] mainOff_add2_rep_bits_out,
    input [9:0] mainOff_add2_rep_tag,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire mainComp_mainOff_add2_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add1_rep_ready;
  wire[9:0] mainComp_mainOff_add1_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add1_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add1_req_bits_in1;
  wire[63:0] mainComp_mainOff_add1_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign mainOff_add2_rep_ready = mainComp_mainOff_add2_rep_ready;
  assign mainOff_add2_req_tag = mainComp_mainOff_add2_req_tag;
  assign mainOff_add2_req_valid = mainComp_mainOff_add2_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_122 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add1_req_ready( offComp_io_in_ready ),
       .mainOff_add1_req_valid( mainComp_mainOff_add1_req_valid ),
       .mainOff_add1_req_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .mainOff_add1_req_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .mainOff_add1_req_tag( mainComp_mainOff_add1_req_tag ),
       .mainOff_add1_rep_ready( mainComp_mainOff_add1_rep_ready ),
       .mainOff_add1_rep_valid( offComp_io_out_valid ),
       .mainOff_add1_rep_bits_out(  ),
       .mainOff_add1_rep_tag( offComp_io_out_tag ),
       .mainOff_add2_req_ready( mainOff_add2_req_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1(  ),
       .mainOff_add2_req_bits_in2(  ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( mainOff_add2_rep_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( mainOff_add2_rep_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_96 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add1_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add1_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add1_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add1_req_tag ),
       .io_out_ready( mainComp_mainOff_add1_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_97(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_97(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_97 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_124(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_sqrt_req_ready,
    output mainOff_sqrt_req_valid,
    output[63:0] mainOff_sqrt_req_bits_in1,
    output[63:0] mainOff_sqrt_req_bits_in2,
    output[9:0] mainOff_sqrt_req_tag,
    output mainOff_sqrt_rep_ready,
    input  mainOff_sqrt_rep_valid,
    input [63:0] mainOff_sqrt_rep_bits_out,
    input [9:0] mainOff_sqrt_rep_tag);

  wire[9:0] mainComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire mainComp_mainOff_sqrt_req_valid;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_add2_rep_ready;
  wire[9:0] mainComp_mainOff_add2_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add2_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_add2_req_bits_in1;
  wire[63:0] mainComp_mainOff_add2_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_sqrt_rep_ready = mainComp_mainOff_sqrt_rep_ready;
  assign mainOff_sqrt_req_tag = mainComp_mainOff_sqrt_req_tag;
  assign mainOff_sqrt_req_valid = mainComp_mainOff_sqrt_req_valid;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_123 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add2_req_ready( offComp_io_in_ready ),
       .mainOff_add2_req_valid( mainComp_mainOff_add2_req_valid ),
       .mainOff_add2_req_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .mainOff_add2_req_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .mainOff_add2_req_tag( mainComp_mainOff_add2_req_tag ),
       .mainOff_add2_rep_ready( mainComp_mainOff_add2_rep_ready ),
       .mainOff_add2_rep_valid( offComp_io_out_valid ),
       .mainOff_add2_rep_bits_out(  ),
       .mainOff_add2_rep_tag( offComp_io_out_tag ),
       .mainOff_sqrt_req_ready( mainOff_sqrt_req_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1(  ),
       .mainOff_sqrt_req_bits_in2(  ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( mainOff_sqrt_rep_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( mainOff_sqrt_rep_tag ));
  FUSynWrapper_97 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add2_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add2_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add2_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add2_req_tag ),
       .io_out_ready( mainComp_mainOff_add2_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_98(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_11;
  reg[4:0] tags_10;
  reg[4:0] tags_9;
  reg[4:0] tags_8;
  reg[4:0] tags_7;
  reg[4:0] tags_6;
  reg[4:0] tags_5;
  reg[4:0] tags_4;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_11;
  reg[0:0] valids_10;
  reg[0:0] valids_9;
  reg[0:0] valids_8;
  reg[0:0] valids_7;
  reg[0:0] valids_6;
  reg[0:0] valids_5;
  reg[0:0] valids_4;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_11};
  assign io_out_valid = valids_11;
  assign io_in_ready = io_out_ready;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_11 <= tags_10;
    end
    if(io_out_ready) begin
      tags_10 <= tags_9;
    end
    if(io_out_ready) begin
      tags_9 <= tags_8;
    end
    if(io_out_ready) begin
      tags_8 <= tags_7;
    end
    if(io_out_ready) begin
      tags_7 <= tags_6;
    end
    if(io_out_ready) begin
      tags_6 <= tags_5;
    end
    if(io_out_ready) begin
      tags_5 <= tags_4;
    end
    if(io_out_ready) begin
      tags_4 <= tags_3;
    end
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_11 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_11 <= valids_10;
    end
    if(reset) begin
      valids_10 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_10 <= valids_9;
    end
    if(reset) begin
      valids_9 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_9 <= valids_8;
    end
    if(reset) begin
      valids_8 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_8 <= valids_7;
    end
    if(reset) begin
      valids_7 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_7 <= valids_6;
    end
    if(reset) begin
      valids_6 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_6 <= valids_5;
    end
    if(reset) begin
      valids_5 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_5 <= valids_4;
    end
    if(reset) begin
      valids_4 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_4 <= valids_3;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_98(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;
  wire tagPipe_io_in_ready;

  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign io_in_ready = tagPipe_io_in_ready;
  assign T1 = 1'h1/* 1*/;
  gPipe_98 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_100_ACMP_dsqrt_4_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_125(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1_x,
    input [63:0] io_in_bits_in1_y,
    input [63:0] io_in_bits_in1_z,
    input [63:0] io_in_bits_in2_x,
    input [63:0] io_in_bits_in2_y,
    input [63:0] io_in_bits_in2_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits_out,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] mainComp_io_out_tag;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_sqrt_rep_ready;
  wire[9:0] mainComp_mainOff_sqrt_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_sqrt_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire mainComp_io_in_ready;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in1;
  wire[63:0] mainComp_mainOff_sqrt_req_bits_in2;

  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_in_ready = mainComp_io_in_ready;
  gOffloadedComponent_124 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_in1_x( io_in_bits_in1_x ),
       .io_in_bits_in1_y( io_in_bits_in1_y ),
       .io_in_bits_in1_z( io_in_bits_in1_z ),
       .io_in_bits_in2_x( io_in_bits_in2_x ),
       .io_in_bits_in2_y( io_in_bits_in2_y ),
       .io_in_bits_in2_z( io_in_bits_in2_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_sqrt_req_ready( offComp_io_in_ready ),
       .mainOff_sqrt_req_valid( mainComp_mainOff_sqrt_req_valid ),
       .mainOff_sqrt_req_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .mainOff_sqrt_req_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .mainOff_sqrt_req_tag( mainComp_mainOff_sqrt_req_tag ),
       .mainOff_sqrt_rep_ready( mainComp_mainOff_sqrt_rep_ready ),
       .mainOff_sqrt_rep_valid( offComp_io_out_valid ),
       .mainOff_sqrt_rep_bits_out(  ),
       .mainOff_sqrt_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_98 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_sqrt_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_sqrt_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_sqrt_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_sqrt_req_tag ),
       .io_out_ready( mainComp_mainOff_sqrt_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gOffloadedComponent_126(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_centeroidMem_req_ready,
    output mainOff_centeroidMem_req_valid,
    output[31:0] mainOff_centeroidMem_req_bits_addr,
    output mainOff_centeroidMem_req_bits_rw,
    output[191:0] mainOff_centeroidMem_req_bits_wData,
    output mainOff_centeroidMem_req_bits_initialize,
    output[9:0] mainOff_centeroidMem_req_tag,
    output mainOff_centeroidMem_rep_ready,
    input  mainOff_centeroidMem_rep_valid,
    input [191:0] mainOff_centeroidMem_rep_bits_rData,
    input [9:0] mainOff_centeroidMem_rep_tag,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire mainComp_mainOff_distanceFU_rep_ready;
  wire mainComp_mainOff_distanceFU_req_valid;
  wire[9:0] mainComp_mainOff_distanceFU_req_tag;
  wire offComp_io_out_valid;
  wire offComp_io_in_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_x;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_x;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_y;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in2_z;
  wire[63:0] mainComp_mainOff_distanceFU_req_bits_in1_z;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign mainOff_centeroidMem_req_tag = mainComp_mainOff_centeroidMem_req_tag;
  assign mainOff_centeroidMem_req_valid = mainComp_mainOff_centeroidMem_req_valid;
  assign mainOff_centeroidMem_rep_ready = mainComp_mainOff_centeroidMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign mainOff_centeroidMem_req_bits_wData = mainComp_mainOff_centeroidMem_req_bits_wData;
  assign mainOff_centeroidMem_req_bits_addr = mainComp_mainOff_centeroidMem_req_bits_addr;
  assign mainOff_centeroidMem_req_bits_rw = mainComp_mainOff_centeroidMem_req_bits_rw;
  KEngine_9 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_distanceFU_req_ready( offComp_io_in_ready ),
       .mainOff_distanceFU_req_valid( mainComp_mainOff_distanceFU_req_valid ),
       .mainOff_distanceFU_req_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .mainOff_distanceFU_req_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .mainOff_distanceFU_req_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .mainOff_distanceFU_req_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .mainOff_distanceFU_req_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .mainOff_distanceFU_req_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .mainOff_distanceFU_req_tag( mainComp_mainOff_distanceFU_req_tag ),
       .mainOff_distanceFU_rep_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .mainOff_distanceFU_rep_valid( offComp_io_out_valid ),
       .mainOff_distanceFU_rep_bits_out(  ),
       .mainOff_distanceFU_rep_tag( offComp_io_out_tag ),
       .mainOff_centeroidMem_req_ready( mainOff_centeroidMem_req_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( mainOff_centeroidMem_rep_valid ),
       .mainOff_centeroidMem_rep_bits_rData( mainOff_centeroidMem_rep_bits_rData ),
       .mainOff_centeroidMem_rep_tag( mainOff_centeroidMem_rep_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  gOffloadedComponent_125 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_distanceFU_req_valid ),
       .io_in_bits_in1_x( mainComp_mainOff_distanceFU_req_bits_in1_x ),
       .io_in_bits_in1_y( mainComp_mainOff_distanceFU_req_bits_in1_y ),
       .io_in_bits_in1_z( mainComp_mainOff_distanceFU_req_bits_in1_z ),
       .io_in_bits_in2_x( mainComp_mainOff_distanceFU_req_bits_in2_x ),
       .io_in_bits_in2_y( mainComp_mainOff_distanceFU_req_bits_in2_y ),
       .io_in_bits_in2_z( mainComp_mainOff_distanceFU_req_bits_in2_z ),
       .io_in_tag( mainComp_mainOff_distanceFU_req_tag ),
       .io_out_ready( mainComp_mainOff_distanceFU_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_out(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_18(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);

  wire[-2:0] T1;
  reg [-2:0] ram [999:0];
  wire[-2:0] T2;
  wire[-2:0] T3;
  wire[-2:0] T6;
  wire[-2:0] T8;
  reg[-2:0] rAddrReg;

  assign io_rData = T0;
  assign T0 = T1;
  assign T1 = ram[T9];
  assign T3 = io_wData;
  assign T4 = T5;
  assign T5 = T6;
  assign T6 = io_rw == T7;
  assign T7 = 1'h1/* 1*/;
  assign T9 = rAddrReg;
  assign T10 = 1'h1/* 1*/;

  always @(posedge clk) begin
    if (T4)
      ram[io_addr] <= T3;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_18(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_18 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_127(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_centeroidMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_centeroidMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_centeroidMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_centeroidMem_req_bits_wData;
  wire[31:0] mainComp_mainOff_centeroidMem_req_bits_addr;
  wire mainComp_mainOff_centeroidMem_req_bits_rw;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_partialAccumulatorMem_req_tag = mainComp_mainOff_partialAccumulatorMem_req_tag;
  assign mainOff_partialAccumulatorMem_req_valid = mainComp_mainOff_partialAccumulatorMem_req_valid;
  assign mainOff_partialAccumulatorMem_rep_ready = mainComp_mainOff_partialAccumulatorMem_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_126 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_centeroidMem_req_ready( offComp_io_in_ready ),
       .mainOff_centeroidMem_req_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .mainOff_centeroidMem_req_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .mainOff_centeroidMem_req_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .mainOff_centeroidMem_req_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .mainOff_centeroidMem_req_bits_initialize(  ),
       .mainOff_centeroidMem_req_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .mainOff_centeroidMem_rep_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .mainOff_centeroidMem_rep_valid( offComp_io_out_valid ),
       .mainOff_centeroidMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_centeroidMem_rep_tag( offComp_io_out_tag ),
       .mainOff_partialAccumulatorMem_req_ready( mainOff_partialAccumulatorMem_req_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( mainOff_partialAccumulatorMem_rep_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( mainOff_partialAccumulatorMem_rep_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_18 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_centeroidMem_req_valid ),
       .io_in_bits_addr( mainComp_mainOff_centeroidMem_req_bits_addr ),
       .io_in_bits_rw( mainComp_mainOff_centeroidMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_centeroidMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_centeroidMem_req_tag ),
       .io_out_ready( mainComp_mainOff_centeroidMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module rawSpMem_19(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [-2:0] io_wData,
    output[-2:0] io_rData);



  always @(posedge clk) begin
  end
endmodule

module spMemComponent_19(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  rawSpMem_19 rspm(.clk(clk), .reset(reset),
       .io_addr(  ),
       .io_rw(  ),
       .io_wData(  ),
       .io_rData(  ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_128(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_127 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr(  ),
       .mainOff_partialAccumulatorMem_req_bits_rw(  ),
       .mainOff_partialAccumulatorMem_req_bits_wData(  ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData(  ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_19 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr(  ),
       .io_in_bits_rw(  ),
       .io_in_bits_wData(  ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_99(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_99(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_99 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_129(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output pcOutN_valid,
    output pcOutN_bits_request,
    output[15:0] pcOutN_bits_moduleId,
    output[7:0] pcOutN_bits_portId,
    output[19:0] pcOutN_bits_pcValue,
    output[3:0] pcOutN_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire mainComp_io_out_valid;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_tag = mainComp_io_out_tag;
  gOffloadedComponent_128 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_99 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gRRDistributor(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_centeroidsFinished,
    output io_out_0_bits_pointsFinished,
    output[15:0] io_out_0_bits_centeroidIndex,
    output[63:0] io_out_0_bits_point_x,
    output[63:0] io_out_0_bits_point_y,
    output[63:0] io_out_0_bits_point_z,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_centeroidsFinished,
    output io_out_1_bits_pointsFinished,
    output[15:0] io_out_1_bits_centeroidIndex,
    output[63:0] io_out_1_bits_point_x,
    output[63:0] io_out_1_bits_point_y,
    output[63:0] io_out_1_bits_point_z,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output io_out_2_bits_centeroidsFinished,
    output io_out_2_bits_pointsFinished,
    output[15:0] io_out_2_bits_centeroidIndex,
    output[63:0] io_out_2_bits_point_x,
    output[63:0] io_out_2_bits_point_y,
    output[63:0] io_out_2_bits_point_z,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output io_out_3_bits_centeroidsFinished,
    output io_out_3_bits_pointsFinished,
    output[15:0] io_out_3_bits_centeroidIndex,
    output[63:0] io_out_3_bits_point_x,
    output[63:0] io_out_3_bits_point_y,
    output[63:0] io_out_3_bits_point_z,
    output[9:0] io_out_3_tag,
    input  io_out_4_ready,
    output io_out_4_valid,
    output io_out_4_bits_centeroidsFinished,
    output io_out_4_bits_pointsFinished,
    output[15:0] io_out_4_bits_centeroidIndex,
    output[63:0] io_out_4_bits_point_x,
    output[63:0] io_out_4_bits_point_y,
    output[63:0] io_out_4_bits_point_z,
    output[9:0] io_out_4_tag,
    input  io_out_5_ready,
    output io_out_5_valid,
    output io_out_5_bits_centeroidsFinished,
    output io_out_5_bits_pointsFinished,
    output[15:0] io_out_5_bits_centeroidIndex,
    output[63:0] io_out_5_bits_point_x,
    output[63:0] io_out_5_bits_point_y,
    output[63:0] io_out_5_bits_point_z,
    output[9:0] io_out_5_tag,
    input  io_out_6_ready,
    output io_out_6_valid,
    output io_out_6_bits_centeroidsFinished,
    output io_out_6_bits_pointsFinished,
    output[15:0] io_out_6_bits_centeroidIndex,
    output[63:0] io_out_6_bits_point_x,
    output[63:0] io_out_6_bits_point_y,
    output[63:0] io_out_6_bits_point_z,
    output[9:0] io_out_6_tag,
    input  io_out_7_ready,
    output io_out_7_valid,
    output io_out_7_bits_centeroidsFinished,
    output io_out_7_bits_pointsFinished,
    output[15:0] io_out_7_bits_centeroidIndex,
    output[63:0] io_out_7_bits_point_x,
    output[63:0] io_out_7_bits_point_y,
    output[63:0] io_out_7_bits_point_z,
    output[9:0] io_out_7_tag,
    input  io_out_8_ready,
    output io_out_8_valid,
    output io_out_8_bits_centeroidsFinished,
    output io_out_8_bits_pointsFinished,
    output[15:0] io_out_8_bits_centeroidIndex,
    output[63:0] io_out_8_bits_point_x,
    output[63:0] io_out_8_bits_point_y,
    output[63:0] io_out_8_bits_point_z,
    output[9:0] io_out_8_tag,
    input  io_out_9_ready,
    output io_out_9_valid,
    output io_out_9_bits_centeroidsFinished,
    output io_out_9_bits_pointsFinished,
    output[15:0] io_out_9_bits_centeroidIndex,
    output[63:0] io_out_9_bits_point_x,
    output[63:0] io_out_9_bits_point_y,
    output[63:0] io_out_9_bits_point_z,
    output[9:0] io_out_9_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    output[3:0] io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  reg[3:0] last_grant;
  wire T43;
  wire[3:0] T44;
  wire[3:0] choose;
  wire[3:0] T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire[3:0] T68;
  wire[3:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[3:0] T74;
  wire T75;
  wire T76;
  wire[3:0] T77;
  wire[3:0] T78;
  wire T79;
  wire T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire T83;
  wire T84;
  wire[3:0] T85;
  wire[3:0] T86;
  wire T87;
  wire T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire T91;
  wire T92;
  wire[3:0] T93;
  wire[3:0] T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  wire T109;
  wire T110;
  wire T111;
  wire[3:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire[3:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire[3:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire[3:0] T124;
  wire T125;
  wire T126;
  wire T127;
  wire[3:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[3:0] T132;
  wire T133;
  wire T134;
  wire[3:0] T135;
  wire T136;
  wire[3:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire[3:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire[3:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire[3:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[3:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire[3:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire[3:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;

  assign io_in_ready = T0;
  assign T0 = T325 || io_out_9_ready;
  assign io_out_9_valid = T1;
  assign T1 = T2 && io_in_valid;
  assign T2 = T314 || T3;
  assign T3 = ! T4;
  assign T4 = T297 || io_out_8_ready;
  assign io_out_8_valid = T5;
  assign T5 = T6 && io_in_valid;
  assign T6 = T287 || T7;
  assign T7 = ! T8;
  assign T8 = T271 || io_out_7_ready;
  assign io_out_7_valid = T9;
  assign T9 = T10 && io_in_valid;
  assign T10 = T261 || T11;
  assign T11 = ! T12;
  assign T12 = T246 || io_out_6_ready;
  assign io_out_6_valid = T13;
  assign T13 = T14 && io_in_valid;
  assign T14 = T237 || T15;
  assign T15 = ! T16;
  assign T16 = T223 || io_out_5_ready;
  assign io_out_5_valid = T17;
  assign T17 = T18 && io_in_valid;
  assign T18 = T215 || T19;
  assign T19 = ! T20;
  assign T20 = T202 || io_out_4_ready;
  assign io_out_4_valid = T21;
  assign T21 = T22 && io_in_valid;
  assign T22 = T195 || T23;
  assign T23 = ! T24;
  assign T24 = T183 || io_out_3_ready;
  assign io_out_3_valid = T25;
  assign T25 = T26 && io_in_valid;
  assign T26 = T177 || T27;
  assign T27 = ! T28;
  assign T28 = T166 || io_out_2_ready;
  assign io_out_2_valid = T29;
  assign T29 = T30 && io_in_valid;
  assign T30 = T161 || T31;
  assign T31 = ! T32;
  assign T32 = T151 || io_out_1_ready;
  assign io_out_1_valid = T33;
  assign T33 = T34 && io_in_valid;
  assign T34 = T147 || T35;
  assign T35 = ! T36;
  assign T36 = T138 || io_out_0_ready;
  assign io_out_0_valid = T37;
  assign T37 = T38 && io_in_valid;
  assign T38 = T136 || T39;
  assign T39 = ! T40;
  assign T40 = T102 || T41;
  assign T41 = io_out_9_ready && T42;
  assign T42 = 4'h9/* 9*/ > last_grant;
  assign T43 = io_in_valid && io_in_ready;
  assign T44 = T43 ? choose : last_grant;
  assign choose = T99 ? T98 : T45;
  assign T45 = T95 ? T94 : T46;
  assign T46 = T91 ? T90 : T47;
  assign T47 = T87 ? T86 : T48;
  assign T48 = T83 ? T82 : T49;
  assign T49 = T79 ? T78 : T50;
  assign T50 = T75 ? T74 : T51;
  assign T51 = T72 ? 4'h8/* 8*/ : T52;
  assign T52 = T70 ? 4'h9/* 9*/ : T53;
  assign T53 = io_out_0_ready ? T69 : T54;
  assign T54 = io_out_1_ready ? T68 : T55;
  assign T55 = io_out_2_ready ? T67 : T56;
  assign T56 = io_out_3_ready ? T66 : T57;
  assign T57 = io_out_4_ready ? T65 : T58;
  assign T58 = io_out_5_ready ? T64 : T59;
  assign T59 = io_out_6_ready ? T63 : T60;
  assign T60 = io_out_7_ready ? T62 : T61;
  assign T61 = io_out_8_ready ? 4'h8/* 8*/ : 4'h9/* 9*/;
  assign T62 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T63 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T64 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T65 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T66 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T67 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T68 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T69 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T70 = io_out_9_ready && T71;
  assign T71 = 4'h9/* 9*/ > last_grant;
  assign T72 = io_out_8_ready && T73;
  assign T73 = 4'h8/* 8*/ > last_grant;
  assign T74 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T75 = io_out_7_ready && T76;
  assign T76 = T77 > last_grant;
  assign T77 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T78 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T79 = io_out_6_ready && T80;
  assign T80 = T81 > last_grant;
  assign T81 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T82 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T83 = io_out_5_ready && T84;
  assign T84 = T85 > last_grant;
  assign T85 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T86 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T87 = io_out_4_ready && T88;
  assign T88 = T89 > last_grant;
  assign T89 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T90 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T91 = io_out_3_ready && T92;
  assign T92 = T93 > last_grant;
  assign T93 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T94 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T95 = io_out_2_ready && T96;
  assign T96 = T97 > last_grant;
  assign T97 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T98 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T99 = io_out_1_ready && T100;
  assign T100 = T101 > last_grant;
  assign T101 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T102 = T105 || T103;
  assign T103 = io_out_8_ready && T104;
  assign T104 = 4'h8/* 8*/ > last_grant;
  assign T105 = T109 || T106;
  assign T106 = io_out_7_ready && T107;
  assign T107 = T108 > last_grant;
  assign T108 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T109 = T113 || T110;
  assign T110 = io_out_6_ready && T111;
  assign T111 = T112 > last_grant;
  assign T112 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T113 = T117 || T114;
  assign T114 = io_out_5_ready && T115;
  assign T115 = T116 > last_grant;
  assign T116 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T117 = T121 || T118;
  assign T118 = io_out_4_ready && T119;
  assign T119 = T120 > last_grant;
  assign T120 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T121 = T125 || T122;
  assign T122 = io_out_3_ready && T123;
  assign T123 = T124 > last_grant;
  assign T124 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T125 = T129 || T126;
  assign T126 = io_out_2_ready && T127;
  assign T127 = T128 > last_grant;
  assign T128 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T129 = T133 || T130;
  assign T130 = io_out_1_ready && T131;
  assign T131 = T132 > last_grant;
  assign T132 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T133 = io_out_0_ready && T134;
  assign T134 = T135 > last_grant;
  assign T135 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T136 = T137 > last_grant;
  assign T137 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign io_out_0_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_0_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T138 = T139 || T41;
  assign T139 = T140 || T103;
  assign T140 = T141 || T106;
  assign T141 = T142 || T110;
  assign T142 = T143 || T114;
  assign T143 = T144 || T118;
  assign T144 = T145 || T122;
  assign T145 = T146 || T126;
  assign T146 = T133 || T130;
  assign T147 = T150 && T148;
  assign T148 = T149 > last_grant;
  assign T149 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T150 = ! T133;
  assign io_out_1_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_1_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T151 = T152 || io_out_0_ready;
  assign T152 = T153 || T41;
  assign T153 = T154 || T103;
  assign T154 = T155 || T106;
  assign T155 = T156 || T110;
  assign T156 = T157 || T114;
  assign T157 = T158 || T118;
  assign T158 = T159 || T122;
  assign T159 = T160 || T126;
  assign T160 = T133 || T130;
  assign T161 = T164 && T162;
  assign T162 = T163 > last_grant;
  assign T163 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T164 = ! T165;
  assign T165 = T133 || T130;
  assign io_out_2_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_2_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T166 = T167 || io_out_1_ready;
  assign T167 = T168 || io_out_0_ready;
  assign T168 = T169 || T41;
  assign T169 = T170 || T103;
  assign T170 = T171 || T106;
  assign T171 = T172 || T110;
  assign T172 = T173 || T114;
  assign T173 = T174 || T118;
  assign T174 = T175 || T122;
  assign T175 = T176 || T126;
  assign T176 = T133 || T130;
  assign T177 = T180 && T178;
  assign T178 = T179 > last_grant;
  assign T179 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T180 = ! T181;
  assign T181 = T182 || T126;
  assign T182 = T133 || T130;
  assign io_out_3_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_3_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T183 = T184 || io_out_2_ready;
  assign T184 = T185 || io_out_1_ready;
  assign T185 = T186 || io_out_0_ready;
  assign T186 = T187 || T41;
  assign T187 = T188 || T103;
  assign T188 = T189 || T106;
  assign T189 = T190 || T110;
  assign T190 = T191 || T114;
  assign T191 = T192 || T118;
  assign T192 = T193 || T122;
  assign T193 = T194 || T126;
  assign T194 = T133 || T130;
  assign T195 = T198 && T196;
  assign T196 = T197 > last_grant;
  assign T197 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T198 = ! T199;
  assign T199 = T200 || T122;
  assign T200 = T201 || T126;
  assign T201 = T133 || T130;
  assign io_out_4_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_4_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T202 = T203 || io_out_3_ready;
  assign T203 = T204 || io_out_2_ready;
  assign T204 = T205 || io_out_1_ready;
  assign T205 = T206 || io_out_0_ready;
  assign T206 = T207 || T41;
  assign T207 = T208 || T103;
  assign T208 = T209 || T106;
  assign T209 = T210 || T110;
  assign T210 = T211 || T114;
  assign T211 = T212 || T118;
  assign T212 = T213 || T122;
  assign T213 = T214 || T126;
  assign T214 = T133 || T130;
  assign T215 = T218 && T216;
  assign T216 = T217 > last_grant;
  assign T217 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T218 = ! T219;
  assign T219 = T220 || T118;
  assign T220 = T221 || T122;
  assign T221 = T222 || T126;
  assign T222 = T133 || T130;
  assign io_out_5_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_5_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T223 = T224 || io_out_4_ready;
  assign T224 = T225 || io_out_3_ready;
  assign T225 = T226 || io_out_2_ready;
  assign T226 = T227 || io_out_1_ready;
  assign T227 = T228 || io_out_0_ready;
  assign T228 = T229 || T41;
  assign T229 = T230 || T103;
  assign T230 = T231 || T106;
  assign T231 = T232 || T110;
  assign T232 = T233 || T114;
  assign T233 = T234 || T118;
  assign T234 = T235 || T122;
  assign T235 = T236 || T126;
  assign T236 = T133 || T130;
  assign T237 = T240 && T238;
  assign T238 = T239 > last_grant;
  assign T239 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T240 = ! T241;
  assign T241 = T242 || T114;
  assign T242 = T243 || T118;
  assign T243 = T244 || T122;
  assign T244 = T245 || T126;
  assign T245 = T133 || T130;
  assign io_out_6_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_6_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T246 = T247 || io_out_5_ready;
  assign T247 = T248 || io_out_4_ready;
  assign T248 = T249 || io_out_3_ready;
  assign T249 = T250 || io_out_2_ready;
  assign T250 = T251 || io_out_1_ready;
  assign T251 = T252 || io_out_0_ready;
  assign T252 = T253 || T41;
  assign T253 = T254 || T103;
  assign T254 = T255 || T106;
  assign T255 = T256 || T110;
  assign T256 = T257 || T114;
  assign T257 = T258 || T118;
  assign T258 = T259 || T122;
  assign T259 = T260 || T126;
  assign T260 = T133 || T130;
  assign T261 = T264 && T262;
  assign T262 = T263 > last_grant;
  assign T263 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T264 = ! T265;
  assign T265 = T266 || T110;
  assign T266 = T267 || T114;
  assign T267 = T268 || T118;
  assign T268 = T269 || T122;
  assign T269 = T270 || T126;
  assign T270 = T133 || T130;
  assign io_out_7_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_7_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T271 = T272 || io_out_6_ready;
  assign T272 = T273 || io_out_5_ready;
  assign T273 = T274 || io_out_4_ready;
  assign T274 = T275 || io_out_3_ready;
  assign T275 = T276 || io_out_2_ready;
  assign T276 = T277 || io_out_1_ready;
  assign T277 = T278 || io_out_0_ready;
  assign T278 = T279 || T41;
  assign T279 = T280 || T103;
  assign T280 = T281 || T106;
  assign T281 = T282 || T110;
  assign T282 = T283 || T114;
  assign T283 = T284 || T118;
  assign T284 = T285 || T122;
  assign T285 = T286 || T126;
  assign T286 = T133 || T130;
  assign T287 = T289 && T288;
  assign T288 = 4'h8/* 8*/ > last_grant;
  assign T289 = ! T290;
  assign T290 = T291 || T106;
  assign T291 = T292 || T110;
  assign T292 = T293 || T114;
  assign T293 = T294 || T118;
  assign T294 = T295 || T122;
  assign T295 = T296 || T126;
  assign T296 = T133 || T130;
  assign io_out_8_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_8_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T297 = T298 || io_out_7_ready;
  assign T298 = T299 || io_out_6_ready;
  assign T299 = T300 || io_out_5_ready;
  assign T300 = T301 || io_out_4_ready;
  assign T301 = T302 || io_out_3_ready;
  assign T302 = T303 || io_out_2_ready;
  assign T303 = T304 || io_out_1_ready;
  assign T304 = T305 || io_out_0_ready;
  assign T305 = T306 || T41;
  assign T306 = T307 || T103;
  assign T307 = T308 || T106;
  assign T308 = T309 || T110;
  assign T309 = T310 || T114;
  assign T310 = T311 || T118;
  assign T311 = T312 || T122;
  assign T312 = T313 || T126;
  assign T313 = T133 || T130;
  assign T314 = T316 && T315;
  assign T315 = 4'h9/* 9*/ > last_grant;
  assign T316 = ! T317;
  assign T317 = T318 || T103;
  assign T318 = T319 || T106;
  assign T319 = T320 || T110;
  assign T320 = T321 || T114;
  assign T321 = T322 || T118;
  assign T322 = T323 || T122;
  assign T323 = T324 || T126;
  assign T324 = T133 || T130;
  assign io_out_9_bits_pointsFinished = io_in_bits_pointsFinished;
  assign io_out_9_bits_centeroidsFinished = io_in_bits_centeroidsFinished;
  assign T325 = T326 || io_out_8_ready;
  assign T326 = T327 || io_out_7_ready;
  assign T327 = T328 || io_out_6_ready;
  assign T328 = T329 || io_out_5_ready;
  assign T329 = T330 || io_out_4_ready;
  assign T330 = T331 || io_out_3_ready;
  assign T331 = T332 || io_out_2_ready;
  assign T332 = io_out_0_ready || io_out_1_ready;
  assign io_out_9_tag = io_in_tag;
  assign io_out_8_tag = io_in_tag;
  assign io_out_7_tag = io_in_tag;
  assign io_out_6_tag = io_in_tag;
  assign io_out_5_tag = io_in_tag;
  assign io_out_4_tag = io_in_tag;
  assign io_out_3_tag = io_in_tag;
  assign io_out_2_tag = io_in_tag;
  assign io_out_1_tag = io_in_tag;
  assign io_out_0_tag = io_in_tag;
  assign io_out_0_bits_point_z = io_in_bits_point_z;
  assign io_out_0_bits_point_y = io_in_bits_point_y;
  assign io_out_0_bits_point_x = io_in_bits_point_x;
  assign io_out_1_bits_point_z = io_in_bits_point_z;
  assign io_out_1_bits_point_y = io_in_bits_point_y;
  assign io_out_1_bits_point_x = io_in_bits_point_x;
  assign io_out_2_bits_point_z = io_in_bits_point_z;
  assign io_out_2_bits_point_y = io_in_bits_point_y;
  assign io_out_2_bits_point_x = io_in_bits_point_x;
  assign io_out_3_bits_point_z = io_in_bits_point_z;
  assign io_out_3_bits_point_y = io_in_bits_point_y;
  assign io_out_3_bits_point_x = io_in_bits_point_x;
  assign io_out_4_bits_point_z = io_in_bits_point_z;
  assign io_out_4_bits_point_y = io_in_bits_point_y;
  assign io_out_4_bits_point_x = io_in_bits_point_x;
  assign io_out_5_bits_point_z = io_in_bits_point_z;
  assign io_out_5_bits_point_y = io_in_bits_point_y;
  assign io_out_5_bits_point_x = io_in_bits_point_x;
  assign io_out_6_bits_point_z = io_in_bits_point_z;
  assign io_out_6_bits_point_y = io_in_bits_point_y;
  assign io_out_6_bits_point_x = io_in_bits_point_x;
  assign io_out_7_bits_point_z = io_in_bits_point_z;
  assign io_out_7_bits_point_y = io_in_bits_point_y;
  assign io_out_7_bits_point_x = io_in_bits_point_x;
  assign io_out_8_bits_point_z = io_in_bits_point_z;
  assign io_out_8_bits_point_y = io_in_bits_point_y;
  assign io_out_8_bits_point_x = io_in_bits_point_x;
  assign io_out_9_bits_point_z = io_in_bits_point_z;
  assign io_out_9_bits_point_y = io_in_bits_point_y;
  assign io_out_9_bits_point_x = io_in_bits_point_x;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 4'h0/* 0*/;
    end else if(T43) begin
      last_grant <= T44;
    end
  end
endmodule

module RRDistributorComponent(input clk, input reset,
    input  io_out_0_ready,
    output io_out_0_valid,
    output io_out_0_bits_centeroidsFinished,
    output io_out_0_bits_pointsFinished,
    output[15:0] io_out_0_bits_centeroidIndex,
    output[63:0] io_out_0_bits_point_x,
    output[63:0] io_out_0_bits_point_y,
    output[63:0] io_out_0_bits_point_z,
    output[9:0] io_out_0_tag,
    input  io_out_1_ready,
    output io_out_1_valid,
    output io_out_1_bits_centeroidsFinished,
    output io_out_1_bits_pointsFinished,
    output[15:0] io_out_1_bits_centeroidIndex,
    output[63:0] io_out_1_bits_point_x,
    output[63:0] io_out_1_bits_point_y,
    output[63:0] io_out_1_bits_point_z,
    output[9:0] io_out_1_tag,
    input  io_out_2_ready,
    output io_out_2_valid,
    output io_out_2_bits_centeroidsFinished,
    output io_out_2_bits_pointsFinished,
    output[15:0] io_out_2_bits_centeroidIndex,
    output[63:0] io_out_2_bits_point_x,
    output[63:0] io_out_2_bits_point_y,
    output[63:0] io_out_2_bits_point_z,
    output[9:0] io_out_2_tag,
    input  io_out_3_ready,
    output io_out_3_valid,
    output io_out_3_bits_centeroidsFinished,
    output io_out_3_bits_pointsFinished,
    output[15:0] io_out_3_bits_centeroidIndex,
    output[63:0] io_out_3_bits_point_x,
    output[63:0] io_out_3_bits_point_y,
    output[63:0] io_out_3_bits_point_z,
    output[9:0] io_out_3_tag,
    input  io_out_4_ready,
    output io_out_4_valid,
    output io_out_4_bits_centeroidsFinished,
    output io_out_4_bits_pointsFinished,
    output[15:0] io_out_4_bits_centeroidIndex,
    output[63:0] io_out_4_bits_point_x,
    output[63:0] io_out_4_bits_point_y,
    output[63:0] io_out_4_bits_point_z,
    output[9:0] io_out_4_tag,
    input  io_out_5_ready,
    output io_out_5_valid,
    output io_out_5_bits_centeroidsFinished,
    output io_out_5_bits_pointsFinished,
    output[15:0] io_out_5_bits_centeroidIndex,
    output[63:0] io_out_5_bits_point_x,
    output[63:0] io_out_5_bits_point_y,
    output[63:0] io_out_5_bits_point_z,
    output[9:0] io_out_5_tag,
    input  io_out_6_ready,
    output io_out_6_valid,
    output io_out_6_bits_centeroidsFinished,
    output io_out_6_bits_pointsFinished,
    output[15:0] io_out_6_bits_centeroidIndex,
    output[63:0] io_out_6_bits_point_x,
    output[63:0] io_out_6_bits_point_y,
    output[63:0] io_out_6_bits_point_z,
    output[9:0] io_out_6_tag,
    input  io_out_7_ready,
    output io_out_7_valid,
    output io_out_7_bits_centeroidsFinished,
    output io_out_7_bits_pointsFinished,
    output[15:0] io_out_7_bits_centeroidIndex,
    output[63:0] io_out_7_bits_point_x,
    output[63:0] io_out_7_bits_point_y,
    output[63:0] io_out_7_bits_point_z,
    output[9:0] io_out_7_tag,
    input  io_out_8_ready,
    output io_out_8_valid,
    output io_out_8_bits_centeroidsFinished,
    output io_out_8_bits_pointsFinished,
    output[15:0] io_out_8_bits_centeroidIndex,
    output[63:0] io_out_8_bits_point_x,
    output[63:0] io_out_8_bits_point_y,
    output[63:0] io_out_8_bits_point_z,
    output[9:0] io_out_8_tag,
    input  io_out_9_ready,
    output io_out_9_valid,
    output io_out_9_bits_centeroidsFinished,
    output io_out_9_bits_pointsFinished,
    output[15:0] io_out_9_bits_centeroidIndex,
    output[63:0] io_out_9_bits_point_x,
    output[63:0] io_out_9_bits_point_y,
    output[63:0] io_out_9_bits_point_z,
    output[9:0] io_out_9_tag,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    output[3:0] io_chosen);

  wire rrDist_io_in_ready;
  wire rrDist_io_out_9_valid;
  wire rrDist_io_out_8_valid;
  wire rrDist_io_out_7_valid;
  wire rrDist_io_out_6_valid;
  wire rrDist_io_out_5_valid;
  wire rrDist_io_out_4_valid;
  wire rrDist_io_out_3_valid;
  wire rrDist_io_out_2_valid;
  wire rrDist_io_out_1_valid;
  wire rrDist_io_out_0_valid;
  wire rrDist_io_out_0_bits_pointsFinished;
  wire rrDist_io_out_0_bits_centeroidsFinished;
  wire rrDist_io_out_1_bits_pointsFinished;
  wire rrDist_io_out_1_bits_centeroidsFinished;
  wire rrDist_io_out_2_bits_pointsFinished;
  wire rrDist_io_out_2_bits_centeroidsFinished;
  wire rrDist_io_out_3_bits_pointsFinished;
  wire rrDist_io_out_3_bits_centeroidsFinished;
  wire rrDist_io_out_4_bits_pointsFinished;
  wire rrDist_io_out_4_bits_centeroidsFinished;
  wire rrDist_io_out_5_bits_pointsFinished;
  wire rrDist_io_out_5_bits_centeroidsFinished;
  wire rrDist_io_out_6_bits_pointsFinished;
  wire rrDist_io_out_6_bits_centeroidsFinished;
  wire rrDist_io_out_7_bits_pointsFinished;
  wire rrDist_io_out_7_bits_centeroidsFinished;
  wire rrDist_io_out_8_bits_pointsFinished;
  wire rrDist_io_out_8_bits_centeroidsFinished;
  wire rrDist_io_out_9_bits_pointsFinished;
  wire rrDist_io_out_9_bits_centeroidsFinished;
  wire[9:0] rrDist_io_out_9_tag;
  wire[9:0] rrDist_io_out_8_tag;
  wire[9:0] rrDist_io_out_7_tag;
  wire[9:0] rrDist_io_out_6_tag;
  wire[9:0] rrDist_io_out_5_tag;
  wire[9:0] rrDist_io_out_4_tag;
  wire[9:0] rrDist_io_out_3_tag;
  wire[9:0] rrDist_io_out_2_tag;
  wire[9:0] rrDist_io_out_1_tag;
  wire[9:0] rrDist_io_out_0_tag;
  wire[63:0] rrDist_io_out_0_bits_point_z;
  wire[63:0] rrDist_io_out_0_bits_point_y;
  wire[63:0] rrDist_io_out_0_bits_point_x;
  wire[63:0] rrDist_io_out_1_bits_point_z;
  wire[63:0] rrDist_io_out_1_bits_point_y;
  wire[63:0] rrDist_io_out_1_bits_point_x;
  wire[63:0] rrDist_io_out_2_bits_point_z;
  wire[63:0] rrDist_io_out_2_bits_point_y;
  wire[63:0] rrDist_io_out_2_bits_point_x;
  wire[63:0] rrDist_io_out_3_bits_point_z;
  wire[63:0] rrDist_io_out_3_bits_point_y;
  wire[63:0] rrDist_io_out_3_bits_point_x;
  wire[63:0] rrDist_io_out_4_bits_point_z;
  wire[63:0] rrDist_io_out_4_bits_point_y;
  wire[63:0] rrDist_io_out_4_bits_point_x;
  wire[63:0] rrDist_io_out_5_bits_point_z;
  wire[63:0] rrDist_io_out_5_bits_point_y;
  wire[63:0] rrDist_io_out_5_bits_point_x;
  wire[63:0] rrDist_io_out_6_bits_point_z;
  wire[63:0] rrDist_io_out_6_bits_point_y;
  wire[63:0] rrDist_io_out_6_bits_point_x;
  wire[63:0] rrDist_io_out_7_bits_point_z;
  wire[63:0] rrDist_io_out_7_bits_point_y;
  wire[63:0] rrDist_io_out_7_bits_point_x;
  wire[63:0] rrDist_io_out_8_bits_point_z;
  wire[63:0] rrDist_io_out_8_bits_point_y;
  wire[63:0] rrDist_io_out_8_bits_point_x;
  wire[63:0] rrDist_io_out_9_bits_point_z;
  wire[63:0] rrDist_io_out_9_bits_point_y;
  wire[63:0] rrDist_io_out_9_bits_point_x;

  assign io_in_ready = rrDist_io_in_ready;
  assign io_out_9_valid = rrDist_io_out_9_valid;
  assign io_out_8_valid = rrDist_io_out_8_valid;
  assign io_out_7_valid = rrDist_io_out_7_valid;
  assign io_out_6_valid = rrDist_io_out_6_valid;
  assign io_out_5_valid = rrDist_io_out_5_valid;
  assign io_out_4_valid = rrDist_io_out_4_valid;
  assign io_out_3_valid = rrDist_io_out_3_valid;
  assign io_out_2_valid = rrDist_io_out_2_valid;
  assign io_out_1_valid = rrDist_io_out_1_valid;
  assign io_out_0_valid = rrDist_io_out_0_valid;
  assign io_out_0_bits_pointsFinished = rrDist_io_out_0_bits_pointsFinished;
  assign io_out_0_bits_centeroidsFinished = rrDist_io_out_0_bits_centeroidsFinished;
  assign io_out_1_bits_pointsFinished = rrDist_io_out_1_bits_pointsFinished;
  assign io_out_1_bits_centeroidsFinished = rrDist_io_out_1_bits_centeroidsFinished;
  assign io_out_2_bits_pointsFinished = rrDist_io_out_2_bits_pointsFinished;
  assign io_out_2_bits_centeroidsFinished = rrDist_io_out_2_bits_centeroidsFinished;
  assign io_out_3_bits_pointsFinished = rrDist_io_out_3_bits_pointsFinished;
  assign io_out_3_bits_centeroidsFinished = rrDist_io_out_3_bits_centeroidsFinished;
  assign io_out_4_bits_pointsFinished = rrDist_io_out_4_bits_pointsFinished;
  assign io_out_4_bits_centeroidsFinished = rrDist_io_out_4_bits_centeroidsFinished;
  assign io_out_5_bits_pointsFinished = rrDist_io_out_5_bits_pointsFinished;
  assign io_out_5_bits_centeroidsFinished = rrDist_io_out_5_bits_centeroidsFinished;
  assign io_out_6_bits_pointsFinished = rrDist_io_out_6_bits_pointsFinished;
  assign io_out_6_bits_centeroidsFinished = rrDist_io_out_6_bits_centeroidsFinished;
  assign io_out_7_bits_pointsFinished = rrDist_io_out_7_bits_pointsFinished;
  assign io_out_7_bits_centeroidsFinished = rrDist_io_out_7_bits_centeroidsFinished;
  assign io_out_8_bits_pointsFinished = rrDist_io_out_8_bits_pointsFinished;
  assign io_out_8_bits_centeroidsFinished = rrDist_io_out_8_bits_centeroidsFinished;
  assign io_out_9_bits_pointsFinished = rrDist_io_out_9_bits_pointsFinished;
  assign io_out_9_bits_centeroidsFinished = rrDist_io_out_9_bits_centeroidsFinished;
  assign io_out_9_tag = rrDist_io_out_9_tag;
  assign io_out_8_tag = rrDist_io_out_8_tag;
  assign io_out_7_tag = rrDist_io_out_7_tag;
  assign io_out_6_tag = rrDist_io_out_6_tag;
  assign io_out_5_tag = rrDist_io_out_5_tag;
  assign io_out_4_tag = rrDist_io_out_4_tag;
  assign io_out_3_tag = rrDist_io_out_3_tag;
  assign io_out_2_tag = rrDist_io_out_2_tag;
  assign io_out_1_tag = rrDist_io_out_1_tag;
  assign io_out_0_tag = rrDist_io_out_0_tag;
  assign io_out_0_bits_point_z = rrDist_io_out_0_bits_point_z;
  assign io_out_0_bits_point_y = rrDist_io_out_0_bits_point_y;
  assign io_out_0_bits_point_x = rrDist_io_out_0_bits_point_x;
  assign io_out_1_bits_point_z = rrDist_io_out_1_bits_point_z;
  assign io_out_1_bits_point_y = rrDist_io_out_1_bits_point_y;
  assign io_out_1_bits_point_x = rrDist_io_out_1_bits_point_x;
  assign io_out_2_bits_point_z = rrDist_io_out_2_bits_point_z;
  assign io_out_2_bits_point_y = rrDist_io_out_2_bits_point_y;
  assign io_out_2_bits_point_x = rrDist_io_out_2_bits_point_x;
  assign io_out_3_bits_point_z = rrDist_io_out_3_bits_point_z;
  assign io_out_3_bits_point_y = rrDist_io_out_3_bits_point_y;
  assign io_out_3_bits_point_x = rrDist_io_out_3_bits_point_x;
  assign io_out_4_bits_point_z = rrDist_io_out_4_bits_point_z;
  assign io_out_4_bits_point_y = rrDist_io_out_4_bits_point_y;
  assign io_out_4_bits_point_x = rrDist_io_out_4_bits_point_x;
  assign io_out_5_bits_point_z = rrDist_io_out_5_bits_point_z;
  assign io_out_5_bits_point_y = rrDist_io_out_5_bits_point_y;
  assign io_out_5_bits_point_x = rrDist_io_out_5_bits_point_x;
  assign io_out_6_bits_point_z = rrDist_io_out_6_bits_point_z;
  assign io_out_6_bits_point_y = rrDist_io_out_6_bits_point_y;
  assign io_out_6_bits_point_x = rrDist_io_out_6_bits_point_x;
  assign io_out_7_bits_point_z = rrDist_io_out_7_bits_point_z;
  assign io_out_7_bits_point_y = rrDist_io_out_7_bits_point_y;
  assign io_out_7_bits_point_x = rrDist_io_out_7_bits_point_x;
  assign io_out_8_bits_point_z = rrDist_io_out_8_bits_point_z;
  assign io_out_8_bits_point_y = rrDist_io_out_8_bits_point_y;
  assign io_out_8_bits_point_x = rrDist_io_out_8_bits_point_x;
  assign io_out_9_bits_point_z = rrDist_io_out_9_bits_point_z;
  assign io_out_9_bits_point_y = rrDist_io_out_9_bits_point_y;
  assign io_out_9_bits_point_x = rrDist_io_out_9_bits_point_x;
  gRRDistributor rrDist(.clk(clk), .reset(reset),
       .io_out_0_ready( io_out_0_ready ),
       .io_out_0_valid( rrDist_io_out_0_valid ),
       .io_out_0_bits_centeroidsFinished( rrDist_io_out_0_bits_centeroidsFinished ),
       .io_out_0_bits_pointsFinished( rrDist_io_out_0_bits_pointsFinished ),
       .io_out_0_bits_centeroidIndex(  ),
       .io_out_0_bits_point_x( rrDist_io_out_0_bits_point_x ),
       .io_out_0_bits_point_y( rrDist_io_out_0_bits_point_y ),
       .io_out_0_bits_point_z( rrDist_io_out_0_bits_point_z ),
       .io_out_0_tag( rrDist_io_out_0_tag ),
       .io_out_1_ready( io_out_1_ready ),
       .io_out_1_valid( rrDist_io_out_1_valid ),
       .io_out_1_bits_centeroidsFinished( rrDist_io_out_1_bits_centeroidsFinished ),
       .io_out_1_bits_pointsFinished( rrDist_io_out_1_bits_pointsFinished ),
       .io_out_1_bits_centeroidIndex(  ),
       .io_out_1_bits_point_x( rrDist_io_out_1_bits_point_x ),
       .io_out_1_bits_point_y( rrDist_io_out_1_bits_point_y ),
       .io_out_1_bits_point_z( rrDist_io_out_1_bits_point_z ),
       .io_out_1_tag( rrDist_io_out_1_tag ),
       .io_out_2_ready( io_out_2_ready ),
       .io_out_2_valid( rrDist_io_out_2_valid ),
       .io_out_2_bits_centeroidsFinished( rrDist_io_out_2_bits_centeroidsFinished ),
       .io_out_2_bits_pointsFinished( rrDist_io_out_2_bits_pointsFinished ),
       .io_out_2_bits_centeroidIndex(  ),
       .io_out_2_bits_point_x( rrDist_io_out_2_bits_point_x ),
       .io_out_2_bits_point_y( rrDist_io_out_2_bits_point_y ),
       .io_out_2_bits_point_z( rrDist_io_out_2_bits_point_z ),
       .io_out_2_tag( rrDist_io_out_2_tag ),
       .io_out_3_ready( io_out_3_ready ),
       .io_out_3_valid( rrDist_io_out_3_valid ),
       .io_out_3_bits_centeroidsFinished( rrDist_io_out_3_bits_centeroidsFinished ),
       .io_out_3_bits_pointsFinished( rrDist_io_out_3_bits_pointsFinished ),
       .io_out_3_bits_centeroidIndex(  ),
       .io_out_3_bits_point_x( rrDist_io_out_3_bits_point_x ),
       .io_out_3_bits_point_y( rrDist_io_out_3_bits_point_y ),
       .io_out_3_bits_point_z( rrDist_io_out_3_bits_point_z ),
       .io_out_3_tag( rrDist_io_out_3_tag ),
       .io_out_4_ready( io_out_4_ready ),
       .io_out_4_valid( rrDist_io_out_4_valid ),
       .io_out_4_bits_centeroidsFinished( rrDist_io_out_4_bits_centeroidsFinished ),
       .io_out_4_bits_pointsFinished( rrDist_io_out_4_bits_pointsFinished ),
       .io_out_4_bits_centeroidIndex(  ),
       .io_out_4_bits_point_x( rrDist_io_out_4_bits_point_x ),
       .io_out_4_bits_point_y( rrDist_io_out_4_bits_point_y ),
       .io_out_4_bits_point_z( rrDist_io_out_4_bits_point_z ),
       .io_out_4_tag( rrDist_io_out_4_tag ),
       .io_out_5_ready( io_out_5_ready ),
       .io_out_5_valid( rrDist_io_out_5_valid ),
       .io_out_5_bits_centeroidsFinished( rrDist_io_out_5_bits_centeroidsFinished ),
       .io_out_5_bits_pointsFinished( rrDist_io_out_5_bits_pointsFinished ),
       .io_out_5_bits_centeroidIndex(  ),
       .io_out_5_bits_point_x( rrDist_io_out_5_bits_point_x ),
       .io_out_5_bits_point_y( rrDist_io_out_5_bits_point_y ),
       .io_out_5_bits_point_z( rrDist_io_out_5_bits_point_z ),
       .io_out_5_tag( rrDist_io_out_5_tag ),
       .io_out_6_ready( io_out_6_ready ),
       .io_out_6_valid( rrDist_io_out_6_valid ),
       .io_out_6_bits_centeroidsFinished( rrDist_io_out_6_bits_centeroidsFinished ),
       .io_out_6_bits_pointsFinished( rrDist_io_out_6_bits_pointsFinished ),
       .io_out_6_bits_centeroidIndex(  ),
       .io_out_6_bits_point_x( rrDist_io_out_6_bits_point_x ),
       .io_out_6_bits_point_y( rrDist_io_out_6_bits_point_y ),
       .io_out_6_bits_point_z( rrDist_io_out_6_bits_point_z ),
       .io_out_6_tag( rrDist_io_out_6_tag ),
       .io_out_7_ready( io_out_7_ready ),
       .io_out_7_valid( rrDist_io_out_7_valid ),
       .io_out_7_bits_centeroidsFinished( rrDist_io_out_7_bits_centeroidsFinished ),
       .io_out_7_bits_pointsFinished( rrDist_io_out_7_bits_pointsFinished ),
       .io_out_7_bits_centeroidIndex(  ),
       .io_out_7_bits_point_x( rrDist_io_out_7_bits_point_x ),
       .io_out_7_bits_point_y( rrDist_io_out_7_bits_point_y ),
       .io_out_7_bits_point_z( rrDist_io_out_7_bits_point_z ),
       .io_out_7_tag( rrDist_io_out_7_tag ),
       .io_out_8_ready( io_out_8_ready ),
       .io_out_8_valid( rrDist_io_out_8_valid ),
       .io_out_8_bits_centeroidsFinished( rrDist_io_out_8_bits_centeroidsFinished ),
       .io_out_8_bits_pointsFinished( rrDist_io_out_8_bits_pointsFinished ),
       .io_out_8_bits_centeroidIndex(  ),
       .io_out_8_bits_point_x( rrDist_io_out_8_bits_point_x ),
       .io_out_8_bits_point_y( rrDist_io_out_8_bits_point_y ),
       .io_out_8_bits_point_z( rrDist_io_out_8_bits_point_z ),
       .io_out_8_tag( rrDist_io_out_8_tag ),
       .io_out_9_ready( io_out_9_ready ),
       .io_out_9_valid( rrDist_io_out_9_valid ),
       .io_out_9_bits_centeroidsFinished( rrDist_io_out_9_bits_centeroidsFinished ),
       .io_out_9_bits_pointsFinished( rrDist_io_out_9_bits_pointsFinished ),
       .io_out_9_bits_centeroidIndex(  ),
       .io_out_9_bits_point_x( rrDist_io_out_9_bits_point_x ),
       .io_out_9_bits_point_y( rrDist_io_out_9_bits_point_y ),
       .io_out_9_bits_point_z( rrDist_io_out_9_bits_point_z ),
       .io_out_9_tag( rrDist_io_out_9_tag ),
       .io_in_ready( rrDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
endmodule

module gRRArbiter(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_centeroidsFinished,
    input  io_in_0_bits_pointsFinished,
    input [15:0] io_in_0_bits_centeroidIndex,
    input [63:0] io_in_0_bits_point_x,
    input [63:0] io_in_0_bits_point_y,
    input [63:0] io_in_0_bits_point_z,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_centeroidsFinished,
    input  io_in_1_bits_pointsFinished,
    input [15:0] io_in_1_bits_centeroidIndex,
    input [63:0] io_in_1_bits_point_x,
    input [63:0] io_in_1_bits_point_y,
    input [63:0] io_in_1_bits_point_z,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_centeroidsFinished,
    input  io_in_2_bits_pointsFinished,
    input [15:0] io_in_2_bits_centeroidIndex,
    input [63:0] io_in_2_bits_point_x,
    input [63:0] io_in_2_bits_point_y,
    input [63:0] io_in_2_bits_point_z,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_centeroidsFinished,
    input  io_in_3_bits_pointsFinished,
    input [15:0] io_in_3_bits_centeroidIndex,
    input [63:0] io_in_3_bits_point_x,
    input [63:0] io_in_3_bits_point_y,
    input [63:0] io_in_3_bits_point_z,
    input [9:0] io_in_3_tag,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits_centeroidsFinished,
    input  io_in_4_bits_pointsFinished,
    input [15:0] io_in_4_bits_centeroidIndex,
    input [63:0] io_in_4_bits_point_x,
    input [63:0] io_in_4_bits_point_y,
    input [63:0] io_in_4_bits_point_z,
    input [9:0] io_in_4_tag,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits_centeroidsFinished,
    input  io_in_5_bits_pointsFinished,
    input [15:0] io_in_5_bits_centeroidIndex,
    input [63:0] io_in_5_bits_point_x,
    input [63:0] io_in_5_bits_point_y,
    input [63:0] io_in_5_bits_point_z,
    input [9:0] io_in_5_tag,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits_centeroidsFinished,
    input  io_in_6_bits_pointsFinished,
    input [15:0] io_in_6_bits_centeroidIndex,
    input [63:0] io_in_6_bits_point_x,
    input [63:0] io_in_6_bits_point_y,
    input [63:0] io_in_6_bits_point_z,
    input [9:0] io_in_6_tag,
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits_centeroidsFinished,
    input  io_in_7_bits_pointsFinished,
    input [15:0] io_in_7_bits_centeroidIndex,
    input [63:0] io_in_7_bits_point_x,
    input [63:0] io_in_7_bits_point_y,
    input [63:0] io_in_7_bits_point_z,
    input [9:0] io_in_7_tag,
    output io_in_8_ready,
    input  io_in_8_valid,
    input  io_in_8_bits_centeroidsFinished,
    input  io_in_8_bits_pointsFinished,
    input [15:0] io_in_8_bits_centeroidIndex,
    input [63:0] io_in_8_bits_point_x,
    input [63:0] io_in_8_bits_point_y,
    input [63:0] io_in_8_bits_point_z,
    input [9:0] io_in_8_tag,
    output io_in_9_ready,
    input  io_in_9_valid,
    input  io_in_9_bits_centeroidsFinished,
    input  io_in_9_bits_pointsFinished,
    input [15:0] io_in_9_bits_centeroidIndex,
    input [63:0] io_in_9_bits_point_x,
    input [63:0] io_in_9_bits_point_y,
    input [63:0] io_in_9_bits_point_z,
    input [9:0] io_in_9_tag,
    output[3:0] io_chosen);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[15:0] T10;
  wire[15:0] T11;
  wire[15:0] T12;
  wire T13;
  wire[9:0] T14;
  wire[24:0] T15;
  wire[3:0] choose;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[3:0] T36;
  wire[3:0] T37;
  wire[3:0] T38;
  wire[3:0] T39;
  wire[3:0] T40;
  wire T41;
  wire T42;
  reg[3:0] last_grant;
  wire T43;
  wire[3:0] T44;
  wire T45;
  wire T46;
  wire[3:0] T47;
  wire T48;
  wire T49;
  wire[3:0] T50;
  wire[3:0] T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire T56;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire[3:0] T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire T72;
  wire T73;
  wire[3:0] T74;
  wire[15:0] dvec_9_centeroidIndex;
  wire[15:0] T75;
  wire[15:0] T76;
  wire[15:0] T77;
  wire T78;
  wire[15:0] dvec_8_centeroidIndex;
  wire[15:0] T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire T82;
  wire[15:0] dvec_7_centeroidIndex;
  wire[15:0] T83;
  wire[15:0] T84;
  wire[15:0] T85;
  wire T86;
  wire[15:0] dvec_6_centeroidIndex;
  wire[15:0] T87;
  wire[15:0] T88;
  wire[15:0] T89;
  wire T90;
  wire[15:0] dvec_5_centeroidIndex;
  wire[15:0] T91;
  wire[15:0] T92;
  wire[15:0] T93;
  wire T94;
  wire[15:0] dvec_4_centeroidIndex;
  wire[15:0] T95;
  wire[15:0] T96;
  wire[15:0] T97;
  wire T98;
  wire[15:0] dvec_3_centeroidIndex;
  wire[15:0] T99;
  wire[15:0] T100;
  wire[15:0] T101;
  wire T102;
  wire[15:0] dvec_2_centeroidIndex;
  wire[15:0] T103;
  wire[15:0] T104;
  wire[15:0] T105;
  wire T106;
  wire[15:0] dvec_1_centeroidIndex;
  wire[15:0] T107;
  wire[15:0] T108;
  wire T109;
  wire[15:0] dvec_0_centeroidIndex;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire[3:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire[3:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire[3:0] T129;
  wire T130;
  wire T131;
  wire T132;
  wire[3:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire[3:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire[3:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire T146;
  wire T147;
  wire[3:0] T148;
  wire T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire[3:0] T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[3:0] T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[3:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire[3:0] T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire[3:0] T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[3:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[3:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire[9:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire T378;
  wire[9:0] T379;
  wire[24:0] T380;
  wire[4:0] tvec_9;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire T385;
  wire[4:0] tvec_8;
  wire[4:0] T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire[4:0] T389;
  wire T390;
  wire[4:0] tvec_7;
  wire[4:0] T391;
  wire[4:0] T392;
  wire[4:0] T393;
  wire[4:0] T394;
  wire T395;
  wire[4:0] tvec_6;
  wire[4:0] T396;
  wire[4:0] T397;
  wire[4:0] T398;
  wire[4:0] T399;
  wire T400;
  wire[4:0] tvec_5;
  wire[4:0] T401;
  wire[4:0] T402;
  wire[4:0] T403;
  wire[4:0] T404;
  wire T405;
  wire[4:0] tvec_4;
  wire[4:0] T406;
  wire[4:0] T407;
  wire[4:0] T408;
  wire[4:0] T409;
  wire T410;
  wire[4:0] tvec_3;
  wire[4:0] T411;
  wire[4:0] T412;
  wire[4:0] T413;
  wire[4:0] T414;
  wire T415;
  wire[4:0] tvec_2;
  wire[4:0] T416;
  wire[4:0] T417;
  wire[4:0] T418;
  wire[4:0] T419;
  wire T420;
  wire[4:0] tvec_1;
  wire[4:0] T421;
  wire[4:0] T422;
  wire[4:0] T423;
  wire T424;
  wire[4:0] tvec_0;
  wire[4:0] T425;

  assign io_in_0_ready = T0;
  assign T0 = T110 && io_out_ready;
  assign io_out_valid = T1;
  assign T1 = T2 || io_in_9_valid;
  assign T2 = T3 || io_in_8_valid;
  assign T3 = T4 || io_in_7_valid;
  assign T4 = T5 || io_in_6_valid;
  assign T5 = T6 || io_in_5_valid;
  assign T6 = T7 || io_in_4_valid;
  assign T7 = T8 || io_in_3_valid;
  assign T8 = T9 || io_in_2_valid;
  assign T9 = io_in_0_valid || io_in_1_valid;
  assign io_out_bits_centeroidIndex = T10;
  assign T10 = T75 | T11;
  assign T11 = dvec_9_centeroidIndex & T12;
  assign T12 = {5'h10/* 16*/{T13}};
  assign T13 = T14[4'h9/* 9*/];
  assign T14 = T15[4'h9/* 9*/:1'h0/* 0*/];
  assign T15 = 10'h1/* 1*/ << choose;
  assign choose = T72 ? T71 : T16;
  assign T16 = T68 ? T67 : T17;
  assign T17 = T64 ? T63 : T18;
  assign T18 = T60 ? T59 : T19;
  assign T19 = T56 ? T55 : T20;
  assign T20 = T52 ? T51 : T21;
  assign T21 = T48 ? T47 : T22;
  assign T22 = T45 ? 4'h8/* 8*/ : T23;
  assign T23 = T41 ? 4'h9/* 9*/ : T24;
  assign T24 = io_in_0_valid ? T40 : T25;
  assign T25 = io_in_1_valid ? T39 : T26;
  assign T26 = io_in_2_valid ? T38 : T27;
  assign T27 = io_in_3_valid ? T37 : T28;
  assign T28 = io_in_4_valid ? T36 : T29;
  assign T29 = io_in_5_valid ? T35 : T30;
  assign T30 = io_in_6_valid ? T34 : T31;
  assign T31 = io_in_7_valid ? T33 : T32;
  assign T32 = io_in_8_valid ? 4'h8/* 8*/ : 4'h9/* 9*/;
  assign T33 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T34 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T35 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T36 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T37 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T38 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T39 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T40 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T41 = io_in_9_valid && T42;
  assign T42 = 4'h9/* 9*/ > last_grant;
  assign T43 = io_out_valid && io_out_ready;
  assign T44 = T43 ? choose : last_grant;
  assign T45 = io_in_8_valid && T46;
  assign T46 = 4'h8/* 8*/ > last_grant;
  assign T47 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T48 = io_in_7_valid && T49;
  assign T49 = T50 > last_grant;
  assign T50 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T51 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T52 = io_in_6_valid && T53;
  assign T53 = T54 > last_grant;
  assign T54 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T55 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T56 = io_in_5_valid && T57;
  assign T57 = T58 > last_grant;
  assign T58 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T59 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T60 = io_in_4_valid && T61;
  assign T61 = T62 > last_grant;
  assign T62 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T63 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T64 = io_in_3_valid && T65;
  assign T65 = T66 > last_grant;
  assign T66 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T67 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T68 = io_in_2_valid && T69;
  assign T69 = T70 > last_grant;
  assign T70 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T71 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T72 = io_in_1_valid && T73;
  assign T73 = T74 > last_grant;
  assign T74 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign dvec_9_centeroidIndex = io_in_9_bits_centeroidIndex;
  assign T75 = T79 | T76;
  assign T76 = dvec_8_centeroidIndex & T77;
  assign T77 = {5'h10/* 16*/{T78}};
  assign T78 = T14[4'h8/* 8*/];
  assign dvec_8_centeroidIndex = io_in_8_bits_centeroidIndex;
  assign T79 = T83 | T80;
  assign T80 = dvec_7_centeroidIndex & T81;
  assign T81 = {5'h10/* 16*/{T82}};
  assign T82 = T14[3'h7/* 7*/];
  assign dvec_7_centeroidIndex = io_in_7_bits_centeroidIndex;
  assign T83 = T87 | T84;
  assign T84 = dvec_6_centeroidIndex & T85;
  assign T85 = {5'h10/* 16*/{T86}};
  assign T86 = T14[3'h6/* 6*/];
  assign dvec_6_centeroidIndex = io_in_6_bits_centeroidIndex;
  assign T87 = T91 | T88;
  assign T88 = dvec_5_centeroidIndex & T89;
  assign T89 = {5'h10/* 16*/{T90}};
  assign T90 = T14[3'h5/* 5*/];
  assign dvec_5_centeroidIndex = io_in_5_bits_centeroidIndex;
  assign T91 = T95 | T92;
  assign T92 = dvec_4_centeroidIndex & T93;
  assign T93 = {5'h10/* 16*/{T94}};
  assign T94 = T14[3'h4/* 4*/];
  assign dvec_4_centeroidIndex = io_in_4_bits_centeroidIndex;
  assign T95 = T99 | T96;
  assign T96 = dvec_3_centeroidIndex & T97;
  assign T97 = {5'h10/* 16*/{T98}};
  assign T98 = T14[2'h3/* 3*/];
  assign dvec_3_centeroidIndex = io_in_3_bits_centeroidIndex;
  assign T99 = T103 | T100;
  assign T100 = dvec_2_centeroidIndex & T101;
  assign T101 = {5'h10/* 16*/{T102}};
  assign T102 = T14[2'h2/* 2*/];
  assign dvec_2_centeroidIndex = io_in_2_bits_centeroidIndex;
  assign T103 = T107 | T104;
  assign T104 = dvec_1_centeroidIndex & T105;
  assign T105 = {5'h10/* 16*/{T106}};
  assign T106 = T14[1'h1/* 1*/];
  assign dvec_1_centeroidIndex = io_in_1_bits_centeroidIndex;
  assign T107 = dvec_0_centeroidIndex & T108;
  assign T108 = {5'h10/* 16*/{T109}};
  assign T109 = T14[1'h0/* 0*/];
  assign dvec_0_centeroidIndex = io_in_0_bits_centeroidIndex;
  assign T110 = T149 || T111;
  assign T111 = ! T112;
  assign T112 = T115 || T113;
  assign T113 = io_in_9_valid && T114;
  assign T114 = 4'h9/* 9*/ > last_grant;
  assign T115 = T118 || T116;
  assign T116 = io_in_8_valid && T117;
  assign T117 = 4'h8/* 8*/ > last_grant;
  assign T118 = T122 || T119;
  assign T119 = io_in_7_valid && T120;
  assign T120 = T121 > last_grant;
  assign T121 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T122 = T126 || T123;
  assign T123 = io_in_6_valid && T124;
  assign T124 = T125 > last_grant;
  assign T125 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T126 = T130 || T127;
  assign T127 = io_in_5_valid && T128;
  assign T128 = T129 > last_grant;
  assign T129 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T130 = T134 || T131;
  assign T131 = io_in_4_valid && T132;
  assign T132 = T133 > last_grant;
  assign T133 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T134 = T138 || T135;
  assign T135 = io_in_3_valid && T136;
  assign T136 = T137 > last_grant;
  assign T137 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T138 = T142 || T139;
  assign T139 = io_in_2_valid && T140;
  assign T140 = T141 > last_grant;
  assign T141 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T142 = T146 || T143;
  assign T143 = io_in_1_valid && T144;
  assign T144 = T145 > last_grant;
  assign T145 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T146 = io_in_0_valid && T147;
  assign T147 = T148 > last_grant;
  assign T148 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign T149 = T150 > last_grant;
  assign T150 = {3'h0/* 0*/, 1'h0/* 0*/};
  assign io_in_1_ready = T151;
  assign T151 = T152 && io_out_ready;
  assign T152 = T164 || T153;
  assign T153 = ! T154;
  assign T154 = T155 || io_in_0_valid;
  assign T155 = T156 || T113;
  assign T156 = T157 || T116;
  assign T157 = T158 || T119;
  assign T158 = T159 || T123;
  assign T159 = T160 || T127;
  assign T160 = T161 || T131;
  assign T161 = T162 || T135;
  assign T162 = T163 || T139;
  assign T163 = T146 || T143;
  assign T164 = T167 && T165;
  assign T165 = T166 > last_grant;
  assign T166 = {3'h0/* 0*/, 1'h1/* 1*/};
  assign T167 = ! T146;
  assign io_in_2_ready = T168;
  assign T168 = T169 && io_out_ready;
  assign T169 = T182 || T170;
  assign T170 = ! T171;
  assign T171 = T172 || io_in_1_valid;
  assign T172 = T173 || io_in_0_valid;
  assign T173 = T174 || T113;
  assign T174 = T175 || T116;
  assign T175 = T176 || T119;
  assign T176 = T177 || T123;
  assign T177 = T178 || T127;
  assign T178 = T179 || T131;
  assign T179 = T180 || T135;
  assign T180 = T181 || T139;
  assign T181 = T146 || T143;
  assign T182 = T185 && T183;
  assign T183 = T184 > last_grant;
  assign T184 = {2'h0/* 0*/, 2'h2/* 2*/};
  assign T185 = ! T186;
  assign T186 = T146 || T143;
  assign io_in_3_ready = T187;
  assign T187 = T188 && io_out_ready;
  assign T188 = T202 || T189;
  assign T189 = ! T190;
  assign T190 = T191 || io_in_2_valid;
  assign T191 = T192 || io_in_1_valid;
  assign T192 = T193 || io_in_0_valid;
  assign T193 = T194 || T113;
  assign T194 = T195 || T116;
  assign T195 = T196 || T119;
  assign T196 = T197 || T123;
  assign T197 = T198 || T127;
  assign T198 = T199 || T131;
  assign T199 = T200 || T135;
  assign T200 = T201 || T139;
  assign T201 = T146 || T143;
  assign T202 = T205 && T203;
  assign T203 = T204 > last_grant;
  assign T204 = {2'h0/* 0*/, 2'h3/* 3*/};
  assign T205 = ! T206;
  assign T206 = T207 || T139;
  assign T207 = T146 || T143;
  assign io_in_4_ready = T208;
  assign T208 = T209 && io_out_ready;
  assign T209 = T224 || T210;
  assign T210 = ! T211;
  assign T211 = T212 || io_in_3_valid;
  assign T212 = T213 || io_in_2_valid;
  assign T213 = T214 || io_in_1_valid;
  assign T214 = T215 || io_in_0_valid;
  assign T215 = T216 || T113;
  assign T216 = T217 || T116;
  assign T217 = T218 || T119;
  assign T218 = T219 || T123;
  assign T219 = T220 || T127;
  assign T220 = T221 || T131;
  assign T221 = T222 || T135;
  assign T222 = T223 || T139;
  assign T223 = T146 || T143;
  assign T224 = T227 && T225;
  assign T225 = T226 > last_grant;
  assign T226 = {1'h0/* 0*/, 3'h4/* 4*/};
  assign T227 = ! T228;
  assign T228 = T229 || T135;
  assign T229 = T230 || T139;
  assign T230 = T146 || T143;
  assign io_in_5_ready = T231;
  assign T231 = T232 && io_out_ready;
  assign T232 = T248 || T233;
  assign T233 = ! T234;
  assign T234 = T235 || io_in_4_valid;
  assign T235 = T236 || io_in_3_valid;
  assign T236 = T237 || io_in_2_valid;
  assign T237 = T238 || io_in_1_valid;
  assign T238 = T239 || io_in_0_valid;
  assign T239 = T240 || T113;
  assign T240 = T241 || T116;
  assign T241 = T242 || T119;
  assign T242 = T243 || T123;
  assign T243 = T244 || T127;
  assign T244 = T245 || T131;
  assign T245 = T246 || T135;
  assign T246 = T247 || T139;
  assign T247 = T146 || T143;
  assign T248 = T251 && T249;
  assign T249 = T250 > last_grant;
  assign T250 = {1'h0/* 0*/, 3'h5/* 5*/};
  assign T251 = ! T252;
  assign T252 = T253 || T131;
  assign T253 = T254 || T135;
  assign T254 = T255 || T139;
  assign T255 = T146 || T143;
  assign io_in_6_ready = T256;
  assign T256 = T257 && io_out_ready;
  assign T257 = T274 || T258;
  assign T258 = ! T259;
  assign T259 = T260 || io_in_5_valid;
  assign T260 = T261 || io_in_4_valid;
  assign T261 = T262 || io_in_3_valid;
  assign T262 = T263 || io_in_2_valid;
  assign T263 = T264 || io_in_1_valid;
  assign T264 = T265 || io_in_0_valid;
  assign T265 = T266 || T113;
  assign T266 = T267 || T116;
  assign T267 = T268 || T119;
  assign T268 = T269 || T123;
  assign T269 = T270 || T127;
  assign T270 = T271 || T131;
  assign T271 = T272 || T135;
  assign T272 = T273 || T139;
  assign T273 = T146 || T143;
  assign T274 = T277 && T275;
  assign T275 = T276 > last_grant;
  assign T276 = {1'h0/* 0*/, 3'h6/* 6*/};
  assign T277 = ! T278;
  assign T278 = T279 || T127;
  assign T279 = T280 || T131;
  assign T280 = T281 || T135;
  assign T281 = T282 || T139;
  assign T282 = T146 || T143;
  assign io_in_7_ready = T283;
  assign T283 = T284 && io_out_ready;
  assign T284 = T302 || T285;
  assign T285 = ! T286;
  assign T286 = T287 || io_in_6_valid;
  assign T287 = T288 || io_in_5_valid;
  assign T288 = T289 || io_in_4_valid;
  assign T289 = T290 || io_in_3_valid;
  assign T290 = T291 || io_in_2_valid;
  assign T291 = T292 || io_in_1_valid;
  assign T292 = T293 || io_in_0_valid;
  assign T293 = T294 || T113;
  assign T294 = T295 || T116;
  assign T295 = T296 || T119;
  assign T296 = T297 || T123;
  assign T297 = T298 || T127;
  assign T298 = T299 || T131;
  assign T299 = T300 || T135;
  assign T300 = T301 || T139;
  assign T301 = T146 || T143;
  assign T302 = T305 && T303;
  assign T303 = T304 > last_grant;
  assign T304 = {1'h0/* 0*/, 3'h7/* 7*/};
  assign T305 = ! T306;
  assign T306 = T307 || T123;
  assign T307 = T308 || T127;
  assign T308 = T309 || T131;
  assign T309 = T310 || T135;
  assign T310 = T311 || T139;
  assign T311 = T146 || T143;
  assign io_in_8_ready = T312;
  assign T312 = T313 && io_out_ready;
  assign T313 = T332 || T314;
  assign T314 = ! T315;
  assign T315 = T316 || io_in_7_valid;
  assign T316 = T317 || io_in_6_valid;
  assign T317 = T318 || io_in_5_valid;
  assign T318 = T319 || io_in_4_valid;
  assign T319 = T320 || io_in_3_valid;
  assign T320 = T321 || io_in_2_valid;
  assign T321 = T322 || io_in_1_valid;
  assign T322 = T323 || io_in_0_valid;
  assign T323 = T324 || T113;
  assign T324 = T325 || T116;
  assign T325 = T326 || T119;
  assign T326 = T327 || T123;
  assign T327 = T328 || T127;
  assign T328 = T329 || T131;
  assign T329 = T330 || T135;
  assign T330 = T331 || T139;
  assign T331 = T146 || T143;
  assign T332 = T334 && T333;
  assign T333 = 4'h8/* 8*/ > last_grant;
  assign T334 = ! T335;
  assign T335 = T336 || T119;
  assign T336 = T337 || T123;
  assign T337 = T338 || T127;
  assign T338 = T339 || T131;
  assign T339 = T340 || T135;
  assign T340 = T341 || T139;
  assign T341 = T146 || T143;
  assign io_in_9_ready = T342;
  assign T342 = T343 && io_out_ready;
  assign T343 = T363 || T344;
  assign T344 = ! T345;
  assign T345 = T346 || io_in_8_valid;
  assign T346 = T347 || io_in_7_valid;
  assign T347 = T348 || io_in_6_valid;
  assign T348 = T349 || io_in_5_valid;
  assign T349 = T350 || io_in_4_valid;
  assign T350 = T351 || io_in_3_valid;
  assign T351 = T352 || io_in_2_valid;
  assign T352 = T353 || io_in_1_valid;
  assign T353 = T354 || io_in_0_valid;
  assign T354 = T355 || T113;
  assign T355 = T356 || T116;
  assign T356 = T357 || T119;
  assign T357 = T358 || T123;
  assign T358 = T359 || T127;
  assign T359 = T360 || T131;
  assign T360 = T361 || T135;
  assign T361 = T362 || T139;
  assign T362 = T146 || T143;
  assign T363 = T365 && T364;
  assign T364 = 4'h9/* 9*/ > last_grant;
  assign T365 = ! T366;
  assign T366 = T367 || T116;
  assign T367 = T368 || T119;
  assign T368 = T369 || T123;
  assign T369 = T370 || T127;
  assign T370 = T371 || T131;
  assign T371 = T372 || T135;
  assign T372 = T373 || T139;
  assign T373 = T146 || T143;
  assign io_out_tag = T374;
  assign T374 = {5'h0/* 0*/, T375};
  assign T375 = T382 | T376;
  assign T376 = tvec_9 & T377;
  assign T377 = {3'h5/* 5*/{T378}};
  assign T378 = T379[4'h9/* 9*/];
  assign T379 = T380[4'h9/* 9*/:1'h0/* 0*/];
  assign T380 = 10'h1/* 1*/ << choose;
  assign tvec_9 = T381;
  assign T381 = io_in_9_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T382 = T387 | T383;
  assign T383 = tvec_8 & T384;
  assign T384 = {3'h5/* 5*/{T385}};
  assign T385 = T379[4'h8/* 8*/];
  assign tvec_8 = T386;
  assign T386 = io_in_8_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T387 = T392 | T388;
  assign T388 = tvec_7 & T389;
  assign T389 = {3'h5/* 5*/{T390}};
  assign T390 = T379[3'h7/* 7*/];
  assign tvec_7 = T391;
  assign T391 = io_in_7_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T392 = T397 | T393;
  assign T393 = tvec_6 & T394;
  assign T394 = {3'h5/* 5*/{T395}};
  assign T395 = T379[3'h6/* 6*/];
  assign tvec_6 = T396;
  assign T396 = io_in_6_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T397 = T402 | T398;
  assign T398 = tvec_5 & T399;
  assign T399 = {3'h5/* 5*/{T400}};
  assign T400 = T379[3'h5/* 5*/];
  assign tvec_5 = T401;
  assign T401 = io_in_5_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T402 = T407 | T403;
  assign T403 = tvec_4 & T404;
  assign T404 = {3'h5/* 5*/{T405}};
  assign T405 = T379[3'h4/* 4*/];
  assign tvec_4 = T406;
  assign T406 = io_in_4_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T407 = T412 | T408;
  assign T408 = tvec_3 & T409;
  assign T409 = {3'h5/* 5*/{T410}};
  assign T410 = T379[2'h3/* 3*/];
  assign tvec_3 = T411;
  assign T411 = io_in_3_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T412 = T417 | T413;
  assign T413 = tvec_2 & T414;
  assign T414 = {3'h5/* 5*/{T415}};
  assign T415 = T379[2'h2/* 2*/];
  assign tvec_2 = T416;
  assign T416 = io_in_2_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T417 = T422 | T418;
  assign T418 = tvec_1 & T419;
  assign T419 = {3'h5/* 5*/{T420}};
  assign T420 = T379[1'h1/* 1*/];
  assign tvec_1 = T421;
  assign T421 = io_in_1_tag[3'h4/* 4*/:1'h0/* 0*/];
  assign T422 = tvec_0 & T423;
  assign T423 = {3'h5/* 5*/{T424}};
  assign T424 = T379[1'h0/* 0*/];
  assign tvec_0 = T425;
  assign T425 = io_in_0_tag[3'h4/* 4*/:1'h0/* 0*/];

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 4'h0/* 0*/;
    end else if(T43) begin
      last_grant <= T44;
    end
  end
endmodule

module RRAggregatorComponent(input clk, input reset,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_centeroidsFinished,
    input  io_in_0_bits_pointsFinished,
    input [15:0] io_in_0_bits_centeroidIndex,
    input [63:0] io_in_0_bits_point_x,
    input [63:0] io_in_0_bits_point_y,
    input [63:0] io_in_0_bits_point_z,
    input [9:0] io_in_0_tag,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_centeroidsFinished,
    input  io_in_1_bits_pointsFinished,
    input [15:0] io_in_1_bits_centeroidIndex,
    input [63:0] io_in_1_bits_point_x,
    input [63:0] io_in_1_bits_point_y,
    input [63:0] io_in_1_bits_point_z,
    input [9:0] io_in_1_tag,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_centeroidsFinished,
    input  io_in_2_bits_pointsFinished,
    input [15:0] io_in_2_bits_centeroidIndex,
    input [63:0] io_in_2_bits_point_x,
    input [63:0] io_in_2_bits_point_y,
    input [63:0] io_in_2_bits_point_z,
    input [9:0] io_in_2_tag,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_centeroidsFinished,
    input  io_in_3_bits_pointsFinished,
    input [15:0] io_in_3_bits_centeroidIndex,
    input [63:0] io_in_3_bits_point_x,
    input [63:0] io_in_3_bits_point_y,
    input [63:0] io_in_3_bits_point_z,
    input [9:0] io_in_3_tag,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits_centeroidsFinished,
    input  io_in_4_bits_pointsFinished,
    input [15:0] io_in_4_bits_centeroidIndex,
    input [63:0] io_in_4_bits_point_x,
    input [63:0] io_in_4_bits_point_y,
    input [63:0] io_in_4_bits_point_z,
    input [9:0] io_in_4_tag,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits_centeroidsFinished,
    input  io_in_5_bits_pointsFinished,
    input [15:0] io_in_5_bits_centeroidIndex,
    input [63:0] io_in_5_bits_point_x,
    input [63:0] io_in_5_bits_point_y,
    input [63:0] io_in_5_bits_point_z,
    input [9:0] io_in_5_tag,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits_centeroidsFinished,
    input  io_in_6_bits_pointsFinished,
    input [15:0] io_in_6_bits_centeroidIndex,
    input [63:0] io_in_6_bits_point_x,
    input [63:0] io_in_6_bits_point_y,
    input [63:0] io_in_6_bits_point_z,
    input [9:0] io_in_6_tag,
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits_centeroidsFinished,
    input  io_in_7_bits_pointsFinished,
    input [15:0] io_in_7_bits_centeroidIndex,
    input [63:0] io_in_7_bits_point_x,
    input [63:0] io_in_7_bits_point_y,
    input [63:0] io_in_7_bits_point_z,
    input [9:0] io_in_7_tag,
    output io_in_8_ready,
    input  io_in_8_valid,
    input  io_in_8_bits_centeroidsFinished,
    input  io_in_8_bits_pointsFinished,
    input [15:0] io_in_8_bits_centeroidIndex,
    input [63:0] io_in_8_bits_point_x,
    input [63:0] io_in_8_bits_point_y,
    input [63:0] io_in_8_bits_point_z,
    input [9:0] io_in_8_tag,
    output io_in_9_ready,
    input  io_in_9_valid,
    input  io_in_9_bits_centeroidsFinished,
    input  io_in_9_bits_pointsFinished,
    input [15:0] io_in_9_bits_centeroidIndex,
    input [63:0] io_in_9_bits_point_x,
    input [63:0] io_in_9_bits_point_y,
    input [63:0] io_in_9_bits_point_z,
    input [9:0] io_in_9_tag,
    output[3:0] io_chosen);

  wire rrArb_io_in_0_ready;
  wire rrArb_io_out_valid;
  wire[15:0] rrArb_io_out_bits_centeroidIndex;
  wire rrArb_io_in_1_ready;
  wire rrArb_io_in_2_ready;
  wire rrArb_io_in_3_ready;
  wire rrArb_io_in_4_ready;
  wire rrArb_io_in_5_ready;
  wire rrArb_io_in_6_ready;
  wire rrArb_io_in_7_ready;
  wire rrArb_io_in_8_ready;
  wire rrArb_io_in_9_ready;
  wire[9:0] rrArb_io_out_tag;

  assign io_in_0_ready = rrArb_io_in_0_ready;
  assign io_out_valid = rrArb_io_out_valid;
  assign io_out_bits_centeroidIndex = rrArb_io_out_bits_centeroidIndex;
  assign io_in_1_ready = rrArb_io_in_1_ready;
  assign io_in_2_ready = rrArb_io_in_2_ready;
  assign io_in_3_ready = rrArb_io_in_3_ready;
  assign io_in_4_ready = rrArb_io_in_4_ready;
  assign io_in_5_ready = rrArb_io_in_5_ready;
  assign io_in_6_ready = rrArb_io_in_6_ready;
  assign io_in_7_ready = rrArb_io_in_7_ready;
  assign io_in_8_ready = rrArb_io_in_8_ready;
  assign io_in_9_ready = rrArb_io_in_9_ready;
  assign io_out_tag = rrArb_io_out_tag;
  gRRArbiter rrArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( rrArb_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( rrArb_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( rrArb_io_out_tag ),
       .io_in_0_ready( rrArb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_valid ),
       .io_in_0_bits_centeroidsFinished(  ),
       .io_in_0_bits_pointsFinished(  ),
       .io_in_0_bits_centeroidIndex( io_in_0_bits_centeroidIndex ),
       .io_in_0_bits_point_x(  ),
       .io_in_0_bits_point_y(  ),
       .io_in_0_bits_point_z(  ),
       .io_in_0_tag( io_in_0_tag ),
       .io_in_1_ready( rrArb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_valid ),
       .io_in_1_bits_centeroidsFinished(  ),
       .io_in_1_bits_pointsFinished(  ),
       .io_in_1_bits_centeroidIndex( io_in_1_bits_centeroidIndex ),
       .io_in_1_bits_point_x(  ),
       .io_in_1_bits_point_y(  ),
       .io_in_1_bits_point_z(  ),
       .io_in_1_tag( io_in_1_tag ),
       .io_in_2_ready( rrArb_io_in_2_ready ),
       .io_in_2_valid( io_in_2_valid ),
       .io_in_2_bits_centeroidsFinished(  ),
       .io_in_2_bits_pointsFinished(  ),
       .io_in_2_bits_centeroidIndex( io_in_2_bits_centeroidIndex ),
       .io_in_2_bits_point_x(  ),
       .io_in_2_bits_point_y(  ),
       .io_in_2_bits_point_z(  ),
       .io_in_2_tag( io_in_2_tag ),
       .io_in_3_ready( rrArb_io_in_3_ready ),
       .io_in_3_valid( io_in_3_valid ),
       .io_in_3_bits_centeroidsFinished(  ),
       .io_in_3_bits_pointsFinished(  ),
       .io_in_3_bits_centeroidIndex( io_in_3_bits_centeroidIndex ),
       .io_in_3_bits_point_x(  ),
       .io_in_3_bits_point_y(  ),
       .io_in_3_bits_point_z(  ),
       .io_in_3_tag( io_in_3_tag ),
       .io_in_4_ready( rrArb_io_in_4_ready ),
       .io_in_4_valid( io_in_4_valid ),
       .io_in_4_bits_centeroidsFinished(  ),
       .io_in_4_bits_pointsFinished(  ),
       .io_in_4_bits_centeroidIndex( io_in_4_bits_centeroidIndex ),
       .io_in_4_bits_point_x(  ),
       .io_in_4_bits_point_y(  ),
       .io_in_4_bits_point_z(  ),
       .io_in_4_tag( io_in_4_tag ),
       .io_in_5_ready( rrArb_io_in_5_ready ),
       .io_in_5_valid( io_in_5_valid ),
       .io_in_5_bits_centeroidsFinished(  ),
       .io_in_5_bits_pointsFinished(  ),
       .io_in_5_bits_centeroidIndex( io_in_5_bits_centeroidIndex ),
       .io_in_5_bits_point_x(  ),
       .io_in_5_bits_point_y(  ),
       .io_in_5_bits_point_z(  ),
       .io_in_5_tag( io_in_5_tag ),
       .io_in_6_ready( rrArb_io_in_6_ready ),
       .io_in_6_valid( io_in_6_valid ),
       .io_in_6_bits_centeroidsFinished(  ),
       .io_in_6_bits_pointsFinished(  ),
       .io_in_6_bits_centeroidIndex( io_in_6_bits_centeroidIndex ),
       .io_in_6_bits_point_x(  ),
       .io_in_6_bits_point_y(  ),
       .io_in_6_bits_point_z(  ),
       .io_in_6_tag( io_in_6_tag ),
       .io_in_7_ready( rrArb_io_in_7_ready ),
       .io_in_7_valid( io_in_7_valid ),
       .io_in_7_bits_centeroidsFinished(  ),
       .io_in_7_bits_pointsFinished(  ),
       .io_in_7_bits_centeroidIndex( io_in_7_bits_centeroidIndex ),
       .io_in_7_bits_point_x(  ),
       .io_in_7_bits_point_y(  ),
       .io_in_7_bits_point_z(  ),
       .io_in_7_tag( io_in_7_tag ),
       .io_in_8_ready( rrArb_io_in_8_ready ),
       .io_in_8_valid( io_in_8_valid ),
       .io_in_8_bits_centeroidsFinished(  ),
       .io_in_8_bits_pointsFinished(  ),
       .io_in_8_bits_centeroidIndex( io_in_8_bits_centeroidIndex ),
       .io_in_8_bits_point_x(  ),
       .io_in_8_bits_point_y(  ),
       .io_in_8_bits_point_z(  ),
       .io_in_8_tag( io_in_8_tag ),
       .io_in_9_ready( rrArb_io_in_9_ready ),
       .io_in_9_valid( io_in_9_valid ),
       .io_in_9_bits_centeroidsFinished(  ),
       .io_in_9_bits_pointsFinished(  ),
       .io_in_9_bits_centeroidIndex( io_in_9_bits_centeroidIndex ),
       .io_in_9_bits_point_x(  ),
       .io_in_9_bits_point_y(  ),
       .io_in_9_bits_point_z(  ),
       .io_in_9_tag( io_in_9_tag ),
       .io_chosen(  ));
endmodule

module gReplicatedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire inputDist_io_in_ready;
  wire gOffloadedComponent_9_io_in_ready;
  wire inputDist_io_out_9_valid;
  wire gOffloadedComponent_8_io_in_ready;
  wire inputDist_io_out_8_valid;
  wire gOffloadedComponent_7_io_in_ready;
  wire inputDist_io_out_7_valid;
  wire gOffloadedComponent_6_io_in_ready;
  wire inputDist_io_out_6_valid;
  wire gOffloadedComponent_5_io_in_ready;
  wire inputDist_io_out_5_valid;
  wire gOffloadedComponent_4_io_in_ready;
  wire inputDist_io_out_4_valid;
  wire gOffloadedComponent_3_io_in_ready;
  wire inputDist_io_out_3_valid;
  wire gOffloadedComponent_2_io_in_ready;
  wire inputDist_io_out_2_valid;
  wire gOffloadedComponent_1_io_in_ready;
  wire inputDist_io_out_1_valid;
  wire gOffloadedComponent_io_in_ready;
  wire inputDist_io_out_0_valid;
  wire inputDist_io_out_0_bits_pointsFinished;
  wire inputDist_io_out_0_bits_centeroidsFinished;
  wire outputArb_io_in_0_ready;
  wire outputArb_io_out_valid;
  wire gOffloadedComponent_9_io_out_valid;
  wire gOffloadedComponent_8_io_out_valid;
  wire gOffloadedComponent_7_io_out_valid;
  wire gOffloadedComponent_6_io_out_valid;
  wire gOffloadedComponent_5_io_out_valid;
  wire gOffloadedComponent_4_io_out_valid;
  wire gOffloadedComponent_3_io_out_valid;
  wire gOffloadedComponent_2_io_out_valid;
  wire gOffloadedComponent_1_io_out_valid;
  wire gOffloadedComponent_io_out_valid;
  wire[15:0] outputArb_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_9_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_8_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_7_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_6_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_5_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_4_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_3_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_2_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_1_io_out_bits_centeroidIndex;
  wire[15:0] gOffloadedComponent_io_out_bits_centeroidIndex;
  wire inputDist_io_out_1_bits_pointsFinished;
  wire inputDist_io_out_1_bits_centeroidsFinished;
  wire outputArb_io_in_1_ready;
  wire inputDist_io_out_2_bits_pointsFinished;
  wire inputDist_io_out_2_bits_centeroidsFinished;
  wire outputArb_io_in_2_ready;
  wire inputDist_io_out_3_bits_pointsFinished;
  wire inputDist_io_out_3_bits_centeroidsFinished;
  wire outputArb_io_in_3_ready;
  wire inputDist_io_out_4_bits_pointsFinished;
  wire inputDist_io_out_4_bits_centeroidsFinished;
  wire outputArb_io_in_4_ready;
  wire inputDist_io_out_5_bits_pointsFinished;
  wire inputDist_io_out_5_bits_centeroidsFinished;
  wire outputArb_io_in_5_ready;
  wire inputDist_io_out_6_bits_pointsFinished;
  wire inputDist_io_out_6_bits_centeroidsFinished;
  wire outputArb_io_in_6_ready;
  wire inputDist_io_out_7_bits_pointsFinished;
  wire inputDist_io_out_7_bits_centeroidsFinished;
  wire outputArb_io_in_7_ready;
  wire inputDist_io_out_8_bits_pointsFinished;
  wire inputDist_io_out_8_bits_centeroidsFinished;
  wire outputArb_io_in_8_ready;
  wire inputDist_io_out_9_bits_pointsFinished;
  wire inputDist_io_out_9_bits_centeroidsFinished;
  wire outputArb_io_in_9_ready;
  wire[9:0] outputArb_io_out_tag;
  wire[9:0] gOffloadedComponent_9_io_out_tag;
  wire[9:0] inputDist_io_out_9_tag;
  wire[9:0] gOffloadedComponent_8_io_out_tag;
  wire[9:0] inputDist_io_out_8_tag;
  wire[9:0] gOffloadedComponent_7_io_out_tag;
  wire[9:0] inputDist_io_out_7_tag;
  wire[9:0] gOffloadedComponent_6_io_out_tag;
  wire[9:0] inputDist_io_out_6_tag;
  wire[9:0] gOffloadedComponent_5_io_out_tag;
  wire[9:0] inputDist_io_out_5_tag;
  wire[9:0] gOffloadedComponent_4_io_out_tag;
  wire[9:0] inputDist_io_out_4_tag;
  wire[9:0] gOffloadedComponent_3_io_out_tag;
  wire[9:0] inputDist_io_out_3_tag;
  wire[9:0] gOffloadedComponent_2_io_out_tag;
  wire[9:0] inputDist_io_out_2_tag;
  wire[9:0] gOffloadedComponent_1_io_out_tag;
  wire[9:0] inputDist_io_out_1_tag;
  wire[9:0] gOffloadedComponent_io_out_tag;
  wire[9:0] inputDist_io_out_0_tag;
  wire[63:0] inputDist_io_out_0_bits_point_z;
  wire[63:0] inputDist_io_out_0_bits_point_y;
  wire[63:0] inputDist_io_out_0_bits_point_x;
  wire[63:0] inputDist_io_out_1_bits_point_z;
  wire[63:0] inputDist_io_out_1_bits_point_y;
  wire[63:0] inputDist_io_out_1_bits_point_x;
  wire[63:0] inputDist_io_out_2_bits_point_z;
  wire[63:0] inputDist_io_out_2_bits_point_y;
  wire[63:0] inputDist_io_out_2_bits_point_x;
  wire[63:0] inputDist_io_out_3_bits_point_z;
  wire[63:0] inputDist_io_out_3_bits_point_y;
  wire[63:0] inputDist_io_out_3_bits_point_x;
  wire[63:0] inputDist_io_out_4_bits_point_z;
  wire[63:0] inputDist_io_out_4_bits_point_y;
  wire[63:0] inputDist_io_out_4_bits_point_x;
  wire[63:0] inputDist_io_out_5_bits_point_z;
  wire[63:0] inputDist_io_out_5_bits_point_y;
  wire[63:0] inputDist_io_out_5_bits_point_x;
  wire[63:0] inputDist_io_out_6_bits_point_z;
  wire[63:0] inputDist_io_out_6_bits_point_y;
  wire[63:0] inputDist_io_out_6_bits_point_x;
  wire[63:0] inputDist_io_out_7_bits_point_z;
  wire[63:0] inputDist_io_out_7_bits_point_y;
  wire[63:0] inputDist_io_out_7_bits_point_x;
  wire[63:0] inputDist_io_out_8_bits_point_z;
  wire[63:0] inputDist_io_out_8_bits_point_y;
  wire[63:0] inputDist_io_out_8_bits_point_x;
  wire[63:0] inputDist_io_out_9_bits_point_z;
  wire[63:0] inputDist_io_out_9_bits_point_y;
  wire[63:0] inputDist_io_out_9_bits_point_x;

  assign io_in_ready = inputDist_io_in_ready;
  assign io_out_valid = outputArb_io_out_valid;
  assign io_out_bits_centeroidIndex = outputArb_io_out_bits_centeroidIndex;
  assign io_out_tag = outputArb_io_out_tag;
  gOffloadedComponent_12 gOffloadedComponent(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_io_in_ready ),
       .io_in_valid( inputDist_io_out_0_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_0_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_0_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_0_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_0_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_0_bits_point_z ),
       .io_in_tag( inputDist_io_out_0_tag ),
       .io_out_ready( outputArb_io_in_0_ready ),
       .io_out_valid( gOffloadedComponent_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_io_out_tag ),
       .pcIn0_valid(  ),
       .pcIn0_bits_request(  ),
       .pcIn0_bits_moduleId(  ),
       .pcIn0_bits_portId(  ),
       .pcIn0_bits_pcValue(  ),
       .pcIn0_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_25 gOffloadedComponent_1(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_1_io_in_ready ),
       .io_in_valid( inputDist_io_out_1_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_1_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_1_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_1_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_1_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_1_bits_point_z ),
       .io_in_tag( inputDist_io_out_1_tag ),
       .io_out_ready( outputArb_io_in_1_ready ),
       .io_out_valid( gOffloadedComponent_1_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_1_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_1_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_38 gOffloadedComponent_2(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_2_io_in_ready ),
       .io_in_valid( inputDist_io_out_2_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_2_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_2_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_2_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_2_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_2_bits_point_z ),
       .io_in_tag( inputDist_io_out_2_tag ),
       .io_out_ready( outputArb_io_in_2_ready ),
       .io_out_valid( gOffloadedComponent_2_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_2_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_2_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_51 gOffloadedComponent_3(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_3_io_in_ready ),
       .io_in_valid( inputDist_io_out_3_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_3_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_3_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_3_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_3_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_3_bits_point_z ),
       .io_in_tag( inputDist_io_out_3_tag ),
       .io_out_ready( outputArb_io_in_3_ready ),
       .io_out_valid( gOffloadedComponent_3_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_3_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_3_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_64 gOffloadedComponent_4(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_4_io_in_ready ),
       .io_in_valid( inputDist_io_out_4_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_4_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_4_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_4_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_4_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_4_bits_point_z ),
       .io_in_tag( inputDist_io_out_4_tag ),
       .io_out_ready( outputArb_io_in_4_ready ),
       .io_out_valid( gOffloadedComponent_4_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_4_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_4_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_77 gOffloadedComponent_5(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_5_io_in_ready ),
       .io_in_valid( inputDist_io_out_5_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_5_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_5_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_5_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_5_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_5_bits_point_z ),
       .io_in_tag( inputDist_io_out_5_tag ),
       .io_out_ready( outputArb_io_in_5_ready ),
       .io_out_valid( gOffloadedComponent_5_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_5_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_5_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_90 gOffloadedComponent_6(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_6_io_in_ready ),
       .io_in_valid( inputDist_io_out_6_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_6_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_6_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_6_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_6_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_6_bits_point_z ),
       .io_in_tag( inputDist_io_out_6_tag ),
       .io_out_ready( outputArb_io_in_6_ready ),
       .io_out_valid( gOffloadedComponent_6_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_6_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_6_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_103 gOffloadedComponent_7(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_7_io_in_ready ),
       .io_in_valid( inputDist_io_out_7_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_7_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_7_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_7_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_7_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_7_bits_point_z ),
       .io_in_tag( inputDist_io_out_7_tag ),
       .io_out_ready( outputArb_io_in_7_ready ),
       .io_out_valid( gOffloadedComponent_7_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_7_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_7_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_116 gOffloadedComponent_8(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_8_io_in_ready ),
       .io_in_valid( inputDist_io_out_8_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_8_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_8_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_8_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_8_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_8_bits_point_z ),
       .io_in_tag( inputDist_io_out_8_tag ),
       .io_out_ready( outputArb_io_in_8_ready ),
       .io_out_valid( gOffloadedComponent_8_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_8_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_8_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_129 gOffloadedComponent_9(.clk(clk), .reset(reset),
       .io_in_ready( gOffloadedComponent_9_io_in_ready ),
       .io_in_valid( inputDist_io_out_9_valid ),
       .io_in_bits_centeroidsFinished( inputDist_io_out_9_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( inputDist_io_out_9_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( inputDist_io_out_9_bits_point_x ),
       .io_in_bits_point_y( inputDist_io_out_9_bits_point_y ),
       .io_in_bits_point_z( inputDist_io_out_9_bits_point_z ),
       .io_in_tag( inputDist_io_out_9_tag ),
       .io_out_ready( outputArb_io_in_9_ready ),
       .io_out_valid( gOffloadedComponent_9_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( gOffloadedComponent_9_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( gOffloadedComponent_9_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .pcOutN_valid(  ),
       .pcOutN_bits_request(  ),
       .pcOutN_bits_moduleId(  ),
       .pcOutN_bits_portId(  ),
       .pcOutN_bits_pcValue(  ),
       .pcOutN_bits_pcType(  ));
  RRDistributorComponent inputDist(.clk(clk), .reset(reset),
       .io_out_0_ready( gOffloadedComponent_io_in_ready ),
       .io_out_0_valid( inputDist_io_out_0_valid ),
       .io_out_0_bits_centeroidsFinished( inputDist_io_out_0_bits_centeroidsFinished ),
       .io_out_0_bits_pointsFinished( inputDist_io_out_0_bits_pointsFinished ),
       .io_out_0_bits_centeroidIndex(  ),
       .io_out_0_bits_point_x( inputDist_io_out_0_bits_point_x ),
       .io_out_0_bits_point_y( inputDist_io_out_0_bits_point_y ),
       .io_out_0_bits_point_z( inputDist_io_out_0_bits_point_z ),
       .io_out_0_tag( inputDist_io_out_0_tag ),
       .io_out_1_ready( gOffloadedComponent_1_io_in_ready ),
       .io_out_1_valid( inputDist_io_out_1_valid ),
       .io_out_1_bits_centeroidsFinished( inputDist_io_out_1_bits_centeroidsFinished ),
       .io_out_1_bits_pointsFinished( inputDist_io_out_1_bits_pointsFinished ),
       .io_out_1_bits_centeroidIndex(  ),
       .io_out_1_bits_point_x( inputDist_io_out_1_bits_point_x ),
       .io_out_1_bits_point_y( inputDist_io_out_1_bits_point_y ),
       .io_out_1_bits_point_z( inputDist_io_out_1_bits_point_z ),
       .io_out_1_tag( inputDist_io_out_1_tag ),
       .io_out_2_ready( gOffloadedComponent_2_io_in_ready ),
       .io_out_2_valid( inputDist_io_out_2_valid ),
       .io_out_2_bits_centeroidsFinished( inputDist_io_out_2_bits_centeroidsFinished ),
       .io_out_2_bits_pointsFinished( inputDist_io_out_2_bits_pointsFinished ),
       .io_out_2_bits_centeroidIndex(  ),
       .io_out_2_bits_point_x( inputDist_io_out_2_bits_point_x ),
       .io_out_2_bits_point_y( inputDist_io_out_2_bits_point_y ),
       .io_out_2_bits_point_z( inputDist_io_out_2_bits_point_z ),
       .io_out_2_tag( inputDist_io_out_2_tag ),
       .io_out_3_ready( gOffloadedComponent_3_io_in_ready ),
       .io_out_3_valid( inputDist_io_out_3_valid ),
       .io_out_3_bits_centeroidsFinished( inputDist_io_out_3_bits_centeroidsFinished ),
       .io_out_3_bits_pointsFinished( inputDist_io_out_3_bits_pointsFinished ),
       .io_out_3_bits_centeroidIndex(  ),
       .io_out_3_bits_point_x( inputDist_io_out_3_bits_point_x ),
       .io_out_3_bits_point_y( inputDist_io_out_3_bits_point_y ),
       .io_out_3_bits_point_z( inputDist_io_out_3_bits_point_z ),
       .io_out_3_tag( inputDist_io_out_3_tag ),
       .io_out_4_ready( gOffloadedComponent_4_io_in_ready ),
       .io_out_4_valid( inputDist_io_out_4_valid ),
       .io_out_4_bits_centeroidsFinished( inputDist_io_out_4_bits_centeroidsFinished ),
       .io_out_4_bits_pointsFinished( inputDist_io_out_4_bits_pointsFinished ),
       .io_out_4_bits_centeroidIndex(  ),
       .io_out_4_bits_point_x( inputDist_io_out_4_bits_point_x ),
       .io_out_4_bits_point_y( inputDist_io_out_4_bits_point_y ),
       .io_out_4_bits_point_z( inputDist_io_out_4_bits_point_z ),
       .io_out_4_tag( inputDist_io_out_4_tag ),
       .io_out_5_ready( gOffloadedComponent_5_io_in_ready ),
       .io_out_5_valid( inputDist_io_out_5_valid ),
       .io_out_5_bits_centeroidsFinished( inputDist_io_out_5_bits_centeroidsFinished ),
       .io_out_5_bits_pointsFinished( inputDist_io_out_5_bits_pointsFinished ),
       .io_out_5_bits_centeroidIndex(  ),
       .io_out_5_bits_point_x( inputDist_io_out_5_bits_point_x ),
       .io_out_5_bits_point_y( inputDist_io_out_5_bits_point_y ),
       .io_out_5_bits_point_z( inputDist_io_out_5_bits_point_z ),
       .io_out_5_tag( inputDist_io_out_5_tag ),
       .io_out_6_ready( gOffloadedComponent_6_io_in_ready ),
       .io_out_6_valid( inputDist_io_out_6_valid ),
       .io_out_6_bits_centeroidsFinished( inputDist_io_out_6_bits_centeroidsFinished ),
       .io_out_6_bits_pointsFinished( inputDist_io_out_6_bits_pointsFinished ),
       .io_out_6_bits_centeroidIndex(  ),
       .io_out_6_bits_point_x( inputDist_io_out_6_bits_point_x ),
       .io_out_6_bits_point_y( inputDist_io_out_6_bits_point_y ),
       .io_out_6_bits_point_z( inputDist_io_out_6_bits_point_z ),
       .io_out_6_tag( inputDist_io_out_6_tag ),
       .io_out_7_ready( gOffloadedComponent_7_io_in_ready ),
       .io_out_7_valid( inputDist_io_out_7_valid ),
       .io_out_7_bits_centeroidsFinished( inputDist_io_out_7_bits_centeroidsFinished ),
       .io_out_7_bits_pointsFinished( inputDist_io_out_7_bits_pointsFinished ),
       .io_out_7_bits_centeroidIndex(  ),
       .io_out_7_bits_point_x( inputDist_io_out_7_bits_point_x ),
       .io_out_7_bits_point_y( inputDist_io_out_7_bits_point_y ),
       .io_out_7_bits_point_z( inputDist_io_out_7_bits_point_z ),
       .io_out_7_tag( inputDist_io_out_7_tag ),
       .io_out_8_ready( gOffloadedComponent_8_io_in_ready ),
       .io_out_8_valid( inputDist_io_out_8_valid ),
       .io_out_8_bits_centeroidsFinished( inputDist_io_out_8_bits_centeroidsFinished ),
       .io_out_8_bits_pointsFinished( inputDist_io_out_8_bits_pointsFinished ),
       .io_out_8_bits_centeroidIndex(  ),
       .io_out_8_bits_point_x( inputDist_io_out_8_bits_point_x ),
       .io_out_8_bits_point_y( inputDist_io_out_8_bits_point_y ),
       .io_out_8_bits_point_z( inputDist_io_out_8_bits_point_z ),
       .io_out_8_tag( inputDist_io_out_8_tag ),
       .io_out_9_ready( gOffloadedComponent_9_io_in_ready ),
       .io_out_9_valid( inputDist_io_out_9_valid ),
       .io_out_9_bits_centeroidsFinished( inputDist_io_out_9_bits_centeroidsFinished ),
       .io_out_9_bits_pointsFinished( inputDist_io_out_9_bits_pointsFinished ),
       .io_out_9_bits_centeroidIndex(  ),
       .io_out_9_bits_point_x( inputDist_io_out_9_bits_point_x ),
       .io_out_9_bits_point_y( inputDist_io_out_9_bits_point_y ),
       .io_out_9_bits_point_z( inputDist_io_out_9_bits_point_z ),
       .io_out_9_tag( inputDist_io_out_9_tag ),
       .io_in_ready( inputDist_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_chosen(  ));
  RRAggregatorComponent outputArb(.clk(clk), .reset(reset),
       .io_out_ready( io_out_ready ),
       .io_out_valid( outputArb_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( outputArb_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( outputArb_io_out_tag ),
       .io_in_0_ready( outputArb_io_in_0_ready ),
       .io_in_0_valid( gOffloadedComponent_io_out_valid ),
       .io_in_0_bits_centeroidsFinished(  ),
       .io_in_0_bits_pointsFinished(  ),
       .io_in_0_bits_centeroidIndex( gOffloadedComponent_io_out_bits_centeroidIndex ),
       .io_in_0_bits_point_x(  ),
       .io_in_0_bits_point_y(  ),
       .io_in_0_bits_point_z(  ),
       .io_in_0_tag( gOffloadedComponent_io_out_tag ),
       .io_in_1_ready( outputArb_io_in_1_ready ),
       .io_in_1_valid( gOffloadedComponent_1_io_out_valid ),
       .io_in_1_bits_centeroidsFinished(  ),
       .io_in_1_bits_pointsFinished(  ),
       .io_in_1_bits_centeroidIndex( gOffloadedComponent_1_io_out_bits_centeroidIndex ),
       .io_in_1_bits_point_x(  ),
       .io_in_1_bits_point_y(  ),
       .io_in_1_bits_point_z(  ),
       .io_in_1_tag( gOffloadedComponent_1_io_out_tag ),
       .io_in_2_ready( outputArb_io_in_2_ready ),
       .io_in_2_valid( gOffloadedComponent_2_io_out_valid ),
       .io_in_2_bits_centeroidsFinished(  ),
       .io_in_2_bits_pointsFinished(  ),
       .io_in_2_bits_centeroidIndex( gOffloadedComponent_2_io_out_bits_centeroidIndex ),
       .io_in_2_bits_point_x(  ),
       .io_in_2_bits_point_y(  ),
       .io_in_2_bits_point_z(  ),
       .io_in_2_tag( gOffloadedComponent_2_io_out_tag ),
       .io_in_3_ready( outputArb_io_in_3_ready ),
       .io_in_3_valid( gOffloadedComponent_3_io_out_valid ),
       .io_in_3_bits_centeroidsFinished(  ),
       .io_in_3_bits_pointsFinished(  ),
       .io_in_3_bits_centeroidIndex( gOffloadedComponent_3_io_out_bits_centeroidIndex ),
       .io_in_3_bits_point_x(  ),
       .io_in_3_bits_point_y(  ),
       .io_in_3_bits_point_z(  ),
       .io_in_3_tag( gOffloadedComponent_3_io_out_tag ),
       .io_in_4_ready( outputArb_io_in_4_ready ),
       .io_in_4_valid( gOffloadedComponent_4_io_out_valid ),
       .io_in_4_bits_centeroidsFinished(  ),
       .io_in_4_bits_pointsFinished(  ),
       .io_in_4_bits_centeroidIndex( gOffloadedComponent_4_io_out_bits_centeroidIndex ),
       .io_in_4_bits_point_x(  ),
       .io_in_4_bits_point_y(  ),
       .io_in_4_bits_point_z(  ),
       .io_in_4_tag( gOffloadedComponent_4_io_out_tag ),
       .io_in_5_ready( outputArb_io_in_5_ready ),
       .io_in_5_valid( gOffloadedComponent_5_io_out_valid ),
       .io_in_5_bits_centeroidsFinished(  ),
       .io_in_5_bits_pointsFinished(  ),
       .io_in_5_bits_centeroidIndex( gOffloadedComponent_5_io_out_bits_centeroidIndex ),
       .io_in_5_bits_point_x(  ),
       .io_in_5_bits_point_y(  ),
       .io_in_5_bits_point_z(  ),
       .io_in_5_tag( gOffloadedComponent_5_io_out_tag ),
       .io_in_6_ready( outputArb_io_in_6_ready ),
       .io_in_6_valid( gOffloadedComponent_6_io_out_valid ),
       .io_in_6_bits_centeroidsFinished(  ),
       .io_in_6_bits_pointsFinished(  ),
       .io_in_6_bits_centeroidIndex( gOffloadedComponent_6_io_out_bits_centeroidIndex ),
       .io_in_6_bits_point_x(  ),
       .io_in_6_bits_point_y(  ),
       .io_in_6_bits_point_z(  ),
       .io_in_6_tag( gOffloadedComponent_6_io_out_tag ),
       .io_in_7_ready( outputArb_io_in_7_ready ),
       .io_in_7_valid( gOffloadedComponent_7_io_out_valid ),
       .io_in_7_bits_centeroidsFinished(  ),
       .io_in_7_bits_pointsFinished(  ),
       .io_in_7_bits_centeroidIndex( gOffloadedComponent_7_io_out_bits_centeroidIndex ),
       .io_in_7_bits_point_x(  ),
       .io_in_7_bits_point_y(  ),
       .io_in_7_bits_point_z(  ),
       .io_in_7_tag( gOffloadedComponent_7_io_out_tag ),
       .io_in_8_ready( outputArb_io_in_8_ready ),
       .io_in_8_valid( gOffloadedComponent_8_io_out_valid ),
       .io_in_8_bits_centeroidsFinished(  ),
       .io_in_8_bits_pointsFinished(  ),
       .io_in_8_bits_centeroidIndex( gOffloadedComponent_8_io_out_bits_centeroidIndex ),
       .io_in_8_bits_point_x(  ),
       .io_in_8_bits_point_y(  ),
       .io_in_8_bits_point_z(  ),
       .io_in_8_tag( gOffloadedComponent_8_io_out_tag ),
       .io_in_9_ready( outputArb_io_in_9_ready ),
       .io_in_9_valid( gOffloadedComponent_9_io_out_valid ),
       .io_in_9_bits_centeroidsFinished(  ),
       .io_in_9_bits_pointsFinished(  ),
       .io_in_9_bits_centeroidIndex( gOffloadedComponent_9_io_out_bits_centeroidIndex ),
       .io_in_9_bits_point_x(  ),
       .io_in_9_bits_point_y(  ),
       .io_in_9_bits_point_z(  ),
       .io_in_9_tag( gOffloadedComponent_9_io_out_tag ),
       .io_chosen(  ));
endmodule

module gChainedComponent(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire source_io_in_ready;
  wire sink_io_in_ready;
  wire source_io_out_valid;
  wire source_io_out_bits_pointsFinished;
  wire source_io_out_bits_centeroidsFinished;
  wire sink_io_out_valid;
  wire[15:0] sink_io_out_bits_centeroidIndex;
  wire[9:0] sink_io_out_tag;
  wire[9:0] source_io_out_tag;
  wire[63:0] source_io_out_bits_point_z;
  wire[63:0] source_io_out_bits_point_y;
  wire[63:0] source_io_out_bits_point_x;

  assign io_in_ready = source_io_in_ready;
  assign io_out_valid = sink_io_out_valid;
  assign io_out_bits_centeroidIndex = sink_io_out_bits_centeroidIndex;
  assign io_out_tag = sink_io_out_tag;
  KDistribute source(.clk(clk), .reset(reset),
       .io_in_ready( source_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( sink_io_in_ready ),
       .io_out_valid( source_io_out_valid ),
       .io_out_bits_centeroidsFinished( source_io_out_bits_centeroidsFinished ),
       .io_out_bits_pointsFinished( source_io_out_bits_pointsFinished ),
       .io_out_bits_centeroidIndex(  ),
       .io_out_bits_point_x( source_io_out_bits_point_x ),
       .io_out_bits_point_y( source_io_out_bits_point_y ),
       .io_out_bits_point_z( source_io_out_bits_point_z ),
       .io_out_tag( source_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gReplicatedComponent sink(.clk(clk), .reset(reset),
       .io_in_ready( sink_io_in_ready ),
       .io_in_valid( source_io_out_valid ),
       .io_in_bits_centeroidsFinished( source_io_out_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( source_io_out_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( source_io_out_bits_point_x ),
       .io_in_bits_point_y( source_io_out_bits_point_y ),
       .io_in_bits_point_z( source_io_out_bits_point_z ),
       .io_in_tag( source_io_out_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( sink_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( sink_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x(  ),
       .io_out_bits_point_y(  ),
       .io_out_bits_point_z(  ),
       .io_out_tag( sink_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module RREncode_63(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_64(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module RREncode_65(
    input  io_valid_0,
    output io_chosen,
    input  io_ready);

  wire choose;

  assign io_chosen = choose;
  assign choose = io_valid_0 ? 1'h0/* 0*/ : 1'h1/* 1*/;
endmodule

module KReduce(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_partialAccumulatorMem_req_ready,
    output mainOff_partialAccumulatorMem_req_valid,
    output[31:0] mainOff_partialAccumulatorMem_req_bits_addr,
    output mainOff_partialAccumulatorMem_req_bits_rw,
    output[191:0] mainOff_partialAccumulatorMem_req_bits_wData,
    output mainOff_partialAccumulatorMem_req_bits_initialize,
    output[9:0] mainOff_partialAccumulatorMem_req_tag,
    output mainOff_partialAccumulatorMem_rep_ready,
    input  mainOff_partialAccumulatorMem_rep_valid,
    input [191:0] mainOff_partialAccumulatorMem_rep_bits_rData,
    input [9:0] mainOff_partialAccumulatorMem_rep_tag,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire T0;
  wire sThreadEncoder_io_chosen;
  wire T1;
  wire T2;
  reg[7:0] State_0;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[1:0] T7;
  wire vThreadEncoder_io_chosen;
  wire T8;
  wire AllOffloadsValid_0;
  wire T9;
  wire T10;
  wire T11;
  reg[0:0] addPortHadValidRequest_0;
  wire T12;
  wire T13;
  wire T14;
  wire addPort_req_valid;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[7:0] T19;
  wire[7:0] T20;
  wire[7:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire rThreadEncoder_io_chosen;
  wire T25;
  reg[0:0] subStateTh_0;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire AllOffloadsReady;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg[0:0] addPortHadReadyRequest;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg[0:0] add_ready_received;
  wire T44;
  wire T45;
  wire addPort_req_ready;
  wire addPort_rep_ready;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire partialAccumulatorMemPort_req_valid;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire[7:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[7:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire[7:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  reg[0:0] partialAccumulatorMem_valid_received_0;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[9:0] T72;
  wire[9:0] partialAccumulatorMemPort_rep_tag;
  wire[9:0] partialAccumulatorMemPort_req_tag;
  wire[9:0] T73;
  wire partialAccumulatorMemPort_rep_valid;
  wire T74;
  wire T75;
  wire[4:0] T76;
  wire T77;
  wire T78;
  reg[0:0] partialAccumulatorMemPortHadReadyRequest;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg[0:0] partialAccumulatorMem_ready_received;
  wire T83;
  wire T84;
  wire partialAccumulatorMemPort_req_ready;
  wire partialAccumulatorMemPort_rep_ready;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire[7:0] T90;
  wire T91;
  wire T92;
  wire T93;
  wire[7:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  reg[0:0] add_valid_received_0;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire[9:0] T103;
  wire[9:0] addPort_rep_tag;
  wire[9:0] addPort_req_tag;
  wire[9:0] T104;
  wire addPort_rep_valid;
  wire T105;
  wire T106;
  wire[4:0] T107;
  wire T108;
  wire T109;
  wire[4:0] T110;
  wire T111;
  wire T112;
  wire[4:0] T113;
  wire T114;
  wire T115;
  wire T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  reg[0:0] partialAccumulatorMemPortHadValidRequest_0;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire[4:0] T124;
  wire T125;
  wire T126;
  wire[4:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire[9:0] T131;
  wire T132;
  wire T133;
  wire T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[7:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire[32:0] T144;
  wire[15:0] T145;
  wire[15:0] T146;
  reg[15:0] inputReg_0_centeroidIndex;
  wire T147;
  wire T148;
  wire T149;
  wire[1:0] T150;
  wire T151;
  wire T152;
  wire[15:0] T153;
  wire T154;
  wire T155;
  wire[7:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire[7:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire[7:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire[7:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[7:0] T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[7:0] T191;
  wire[7:0] T192;
  wire[7:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[7:0] T196;
  wire[7:0] T197;
  wire[7:0] T198;
  wire[7:0] T199;
  wire[7:0] T200;
  wire[7:0] T201;
  wire[7:0] T202;
  reg[7:0] EmitReturnState_0;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire[31:0] T208;
  wire[31:0] T209;
  reg[31:0] centeroidIndex_0;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[31:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire T218;
  wire[31:0] T219;
  wire[7:0] T220;
  wire[7:0] T221;
  wire[7:0] T222;
  wire[7:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  wire[7:0] T226;
  wire[7:0] T227;
  wire T228;
  wire[9:0] T229;
  wire[9:0] T230;
  reg[9:0] inputTag_0;
  wire[9:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  reg[0:0] outputReg_0_pointsFinished;
  wire T236;
  wire[15:0] T237;
  wire[15:0] T238;
  reg[15:0] outputReg_0_centeroidIndex;
  wire[15:0] T239;
  wire T240;
  reg[0:0] outputReg_0_centeroidsFinished;
  wire T241;
  wire[63:0] T242;
  wire[63:0] T243;
  reg[63:0] outputReg_0_point_y;
  wire[63:0] T244;
  wire[63:0] T245;
  wire[191:0] T246;
  wire[191:0] T247;
  wire[191:0] T248;
  reg[191:0] pMemOut_0_rData;
  wire T249;
  wire T250;
  wire T251;
  wire[191:0] T252;
  wire[191:0] T253;
  wire[191:0] partialAccumulatorMemPortReplyValue;
  wire[191:0] T254;
  wire[191:0] T255;
  wire[191:0] T256;
  reg[191:0] partialAccumulatorMemPortReplyStorage_0_rData;
  wire T257;
  wire T258;
  wire T259;
  wire[1023:0] T260;
  wire[191:0] T261;
  wire[191:0] partialAccumulatorMemPort_rep_bits_rData;
  wire[191:0] partialAccumulatorMemPort_req_bits_wData;
  wire[191:0] T262;
  wire[225:0] T263;
  wire[225:0] T264;
  wire T265;
  wire[225:0] T266;
  wire[225:0] T267;
  wire T268;
  wire[225:0] T269;
  wire[225:0] T270;
  wire[225:0] T271;
  wire pMemIn3_initialize;
  wire[191:0] pMemIn3_wData;
  wire pMemIn3_rw;
  wire[31:0] pMemIn3_addr;
  wire[31:0] T272;
  wire[31:0] T273;
  wire T274;
  wire T275;
  wire[7:0] T276;
  wire T277;
  wire[191:0] T278;
  wire T279;
  wire[31:0] T280;
  wire[225:0] T281;
  wire pMemIn2_initialize;
  wire[191:0] pMemIn2_wData;
  wire[191:0] T282;
  wire[191:0] T283;
  wire[63:0] T284;
  wire[63:0] T285;
  reg[63:0] memData_0_z;
  wire T286;
  wire[63:0] T287;
  wire[63:0] T288;
  wire[63:0] T289;
  wire[191:0] T290;
  wire[63:0] addOut3_out;
  wire[63:0] T291;
  wire[63:0] addPortReplyValue;
  wire[63:0] T292;
  wire[63:0] T293;
  wire[63:0] T294;
  reg[63:0] addPortReplyStorage_0_out;
  wire T295;
  wire T296;
  wire T297;
  wire[1023:0] T298;
  wire[63:0] T299;
  wire[63:0] addPort_rep_bits_out;
  wire[63:0] T300;
  wire T301;
  wire T302;
  wire[9:0] T303;
  wire[63:0] T304;
  wire[63:0] T305;
  reg[63:0] memData_0_y;
  wire T306;
  wire[63:0] T307;
  wire[63:0] T308;
  wire[63:0] T309;
  wire[63:0] addOut2_out;
  wire[63:0] T310;
  wire[63:0] T311;
  reg[63:0] memData_0_x;
  wire T312;
  wire[63:0] T313;
  wire[63:0] T314;
  wire[63:0] T315;
  wire[63:0] addOut1_out;
  wire pMemIn2_rw;
  wire[31:0] pMemIn2_addr;
  wire[31:0] T316;
  wire[15:0] T317;
  wire[15:0] T318;
  wire T319;
  wire T320;
  wire[7:0] T321;
  wire T322;
  wire[191:0] T323;
  wire T324;
  wire[31:0] T325;
  wire[225:0] T326;
  wire pMemIn1_initialize;
  wire[191:0] pMemIn1_wData;
  wire pMemIn1_rw;
  wire[31:0] pMemIn1_addr;
  wire[31:0] T327;
  wire T328;
  wire T329;
  wire[7:0] T330;
  wire T331;
  wire[31:0] partialAccumulatorMemPort_req_bits_addr;
  wire[31:0] T332;
  wire partialAccumulatorMemPort_req_bits_rw;
  wire T333;
  wire[191:0] T334;
  wire T335;
  wire T336;
  wire[9:0] T337;
  wire T338;
  wire T339;
  wire[63:0] T340;
  wire[63:0] T341;
  reg[63:0] outputReg_0_point_z;
  wire[63:0] T342;
  wire[63:0] T343;
  wire[63:0] T344;
  wire[63:0] T345;
  reg[63:0] outputReg_0_point_x;
  wire[63:0] T346;
  wire[63:0] T347;

  assign io_in_ready = T0;
  assign T0 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T1 = T228 && T2;
  assign T2 = State_0 == 8'h0/* 0*/;
  assign T3 = T139 || T4;
  assign T4 = T133 && T5;
  assign T5 = T6;
  assign T6 = T7[1'h0/* 0*/:1'h0/* 0*/];
  assign T7 = 1'h1/* 1*/ << vThreadEncoder_io_chosen;
  assign T8 = T132 && AllOffloadsValid_0;
  assign AllOffloadsValid_0 = T9;
  assign T9 = T118 && T10;
  assign T10 = T114 || T11;
  assign T11 = ! addPortHadValidRequest_0;
  assign T12 = T111 && T13;
  assign T13 = addPortHadValidRequest_0 || T14;
  assign T14 = T109 && addPort_req_valid;
  assign addPort_req_valid = T15;
  assign T15 = T96 && T16;
  assign T16 = T87 || T17;
  assign T17 = T86 && T18;
  assign T18 = T20 == T19;
  assign T19 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T20 = State_0 & T21;
  assign T21 = {4'h8/* 8*/{T22}};
  assign T22 = T23;
  assign T23 = T24[1'h0/* 0*/:1'h0/* 0*/];
  assign T24 = 1'h1/* 1*/ << rThreadEncoder_io_chosen;
  assign T25 = subStateTh_0 == 1'h0/* 0*/;
  assign T26 = T29 ? 1'h1/* 1*/ : T27;
  assign T27 = T28 ? 1'h0/* 0*/ : subStateTh_0;
  assign T28 = 1'h0/* 0*/ == vThreadEncoder_io_chosen;
  assign T29 = T31 && T30;
  assign T30 = State_0 != 8'hff/* 255*/;
  assign T31 = T33 && T32;
  assign T32 = State_0 != 8'h0/* 0*/;
  assign T33 = AllOffloadsReady && T34;
  assign T34 = 1'h0/* 0*/ == rThreadEncoder_io_chosen;
  assign AllOffloadsReady = T35;
  assign T35 = T47 && T36;
  assign T36 = T43 || T37;
  assign T37 = T39 && T38;
  assign T38 = ! addPort_req_valid;
  assign T39 = ! addPortHadReadyRequest;
  assign T40 = T42 && T41;
  assign T41 = addPortHadReadyRequest || addPort_req_valid;
  assign T42 = ! AllOffloadsReady;
  assign T43 = addPort_req_ready || add_ready_received;
  assign T44 = T46 && T45;
  assign T45 = add_ready_received || addPort_req_ready;
  assign addPort_req_ready = mainOff_add_req_ready;
  assign mainOff_add_rep_ready = addPort_rep_ready;
  assign addPort_rep_ready = 1'h1/* 1*/;
  assign T46 = ! AllOffloadsReady;
  assign T47 = T82 || T48;
  assign T48 = T78 && T49;
  assign T49 = ! partialAccumulatorMemPort_req_valid;
  assign partialAccumulatorMemPort_req_valid = T50;
  assign T50 = T65 && T51;
  assign T51 = T56 || T52;
  assign T52 = T55 && T53;
  assign T53 = T20 == T54;
  assign T54 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T55 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T56 = T61 || T57;
  assign T57 = T60 && T58;
  assign T58 = T20 == T59;
  assign T59 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T60 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T61 = T64 && T62;
  assign T62 = T20 == T63;
  assign T63 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T64 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T65 = T77 && T66;
  assign T66 = ! T67;
  assign T67 = partialAccumulatorMem_valid_received_0 & T22;
  assign T68 = T74 && T69;
  assign T69 = partialAccumulatorMem_valid_received_0 || T70;
  assign T70 = partialAccumulatorMemPort_rep_valid && T71;
  assign T71 = partialAccumulatorMemPort_rep_tag == T72;
  assign T72 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign partialAccumulatorMemPort_rep_tag = mainOff_partialAccumulatorMem_rep_tag;
  assign mainOff_partialAccumulatorMem_req_tag = partialAccumulatorMemPort_req_tag;
  assign partialAccumulatorMemPort_req_tag = T73;
  assign T73 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign partialAccumulatorMemPort_rep_valid = mainOff_partialAccumulatorMem_rep_valid;
  assign mainOff_partialAccumulatorMem_req_valid = partialAccumulatorMemPort_req_valid;
  assign T74 = ! T75;
  assign T75 = T76 == 5'h0/* 0*/;
  assign T76 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T77 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T78 = ! partialAccumulatorMemPortHadReadyRequest;
  assign T79 = T81 && T80;
  assign T80 = partialAccumulatorMemPortHadReadyRequest || partialAccumulatorMemPort_req_valid;
  assign T81 = ! AllOffloadsReady;
  assign T82 = partialAccumulatorMemPort_req_ready || partialAccumulatorMem_ready_received;
  assign T83 = T85 && T84;
  assign T84 = partialAccumulatorMem_ready_received || partialAccumulatorMemPort_req_ready;
  assign partialAccumulatorMemPort_req_ready = mainOff_partialAccumulatorMem_req_ready;
  assign mainOff_partialAccumulatorMem_rep_ready = partialAccumulatorMemPort_rep_ready;
  assign partialAccumulatorMemPort_rep_ready = 1'h1/* 1*/;
  assign T85 = ! AllOffloadsReady;
  assign T86 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T87 = T92 || T88;
  assign T88 = T91 && T89;
  assign T89 = T20 == T90;
  assign T90 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T91 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T92 = T95 && T93;
  assign T93 = T20 == T94;
  assign T94 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T95 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T96 = T108 && T97;
  assign T97 = ! T98;
  assign T98 = add_valid_received_0 & T22;
  assign T99 = T105 && T100;
  assign T100 = add_valid_received_0 || T101;
  assign T101 = addPort_rep_valid && T102;
  assign T102 = addPort_rep_tag == T103;
  assign T103 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign addPort_rep_tag = mainOff_add_rep_tag;
  assign mainOff_add_req_tag = addPort_req_tag;
  assign addPort_req_tag = T104;
  assign T104 = {9'h0/* 0*/, rThreadEncoder_io_chosen};
  assign addPort_rep_valid = mainOff_add_rep_valid;
  assign mainOff_add_req_valid = addPort_req_valid;
  assign T105 = ! T106;
  assign T106 = T107 == 5'h0/* 0*/;
  assign T107 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T108 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T109 = 5'h0/* 0*/ == T110;
  assign T110 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T111 = ! T112;
  assign T112 = T113 == 5'h0/* 0*/;
  assign T113 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T114 = T115 || add_valid_received_0;
  assign T115 = addPort_rep_valid && T116;
  assign T116 = addPort_rep_tag == T117;
  assign T117 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T118 = T128 || T119;
  assign T119 = ! partialAccumulatorMemPortHadValidRequest_0;
  assign T120 = T125 && T121;
  assign T121 = partialAccumulatorMemPortHadValidRequest_0 || T122;
  assign T122 = T123 && partialAccumulatorMemPort_req_valid;
  assign T123 = 5'h0/* 0*/ == T124;
  assign T124 = {4'h0/* 0*/, rThreadEncoder_io_chosen};
  assign T125 = ! T126;
  assign T126 = T127 == 5'h0/* 0*/;
  assign T127 = {4'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T128 = T129 || partialAccumulatorMem_valid_received_0;
  assign T129 = partialAccumulatorMemPort_rep_valid && T130;
  assign T130 = partialAccumulatorMemPort_rep_tag == T131;
  assign T131 = {5'h0/* 0*/, 5'h0/* 0*/};
  assign T132 = subStateTh_0 == 1'h1/* 1*/;
  assign T133 = T138 && T134;
  assign T134 = T136 == T135;
  assign T135 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T136 = State_0 & T137;
  assign T137 = {4'h8/* 8*/{T5}};
  assign T138 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T139 = T158 || T140;
  assign T140 = T141 && T5;
  assign T141 = T154 && T142;
  assign T142 = ! T143;
  assign T143 = T144 == 33'h4/* 4*/;
  assign T144 = {17'h0/* 0*/, T145};
  assign T145 = inputReg_0_centeroidIndex & T146;
  assign T146 = {5'h10/* 16*/{T5}};
  assign T147 = T151 && T148;
  assign T148 = T149;
  assign T149 = T150[1'h0/* 0*/:1'h0/* 0*/];
  assign T150 = 1'h1/* 1*/ << sThreadEncoder_io_chosen;
  assign T151 = T152 && io_in_valid;
  assign T152 = sThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T153 = T147 ? io_in_bits_centeroidIndex : inputReg_0_centeroidIndex;
  assign T154 = T157 && T155;
  assign T155 = T136 == T156;
  assign T156 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T157 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T158 = T161 || T159;
  assign T159 = T160 && T5;
  assign T160 = T154 && T143;
  assign T161 = T167 || T162;
  assign T162 = T163 && T5;
  assign T163 = T166 && T164;
  assign T164 = T136 == T165;
  assign T165 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T166 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T167 = T173 || T168;
  assign T168 = T169 && T5;
  assign T169 = T172 && T170;
  assign T170 = T136 == T171;
  assign T171 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T172 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T173 = T179 || T174;
  assign T174 = T175 && T5;
  assign T175 = T178 && T176;
  assign T176 = T136 == T177;
  assign T177 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T178 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T179 = T185 || T180;
  assign T180 = T181 && T5;
  assign T181 = T184 && T182;
  assign T182 = T136 == T183;
  assign T183 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T184 = vThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T185 = T147 || T186;
  assign T186 = T187 && T22;
  assign T187 = T188 && io_out_ready;
  assign T188 = T190 && T189;
  assign T189 = T20 == 8'hff/* 255*/;
  assign T190 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T191 = T4 ? 8'hff/* 255*/ : T192;
  assign T192 = T140 ? 8'h0/* 0*/ : T193;
  assign T193 = T159 ? T227 : T194;
  assign T194 = T162 ? T226 : T195;
  assign T195 = T168 ? T225 : T196;
  assign T196 = T174 ? T224 : T197;
  assign T197 = T180 ? T223 : T198;
  assign T198 = T186 ? T201 : T199;
  assign T199 = T147 ? T200 : State_0;
  assign T200 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T201 = EmitReturnState_0 & T202;
  assign T202 = {4'h8/* 8*/{T22}};
  assign T203 = T211 || T204;
  assign T204 = T205 && T5;
  assign T205 = T133 && T206;
  assign T206 = ! T207;
  assign T207 = T208 == 32'h5/* 5*/;
  assign T208 = centeroidIndex_0 & T209;
  assign T209 = {6'h20/* 32*/{T5}};
  assign T210 = T213 || T211;
  assign T211 = T212 && T5;
  assign T212 = T133 && T207;
  assign T213 = T214 || T4;
  assign T214 = T147 || T159;
  assign T215 = T211 ? 32'h0/* 0*/ : T216;
  assign T216 = T4 ? T219 : T217;
  assign T217 = T218 ? 32'h0/* 0*/ : centeroidIndex_0;
  assign T218 = T147 || T159;
  assign T219 = T208 + 32'h1/* 1*/;
  assign T220 = T204 ? T222 : T221;
  assign T221 = T211 ? 8'h0/* 0*/ : EmitReturnState_0;
  assign T222 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T223 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign T224 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign T225 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign T226 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T227 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T228 = subStateTh_0 == 1'h0/* 0*/;
  assign io_out_tag = T229;
  assign T229 = inputTag_0 & T230;
  assign T230 = {4'ha/* 10*/{T22}};
  assign T231 = T147 ? io_in_tag : inputTag_0;
  assign io_out_valid = T232;
  assign T232 = T234 && T233;
  assign T233 = T20 == 8'hff/* 255*/;
  assign T234 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign io_out_bits_pointsFinished = T235;
  assign T235 = outputReg_0_pointsFinished & T22;
  assign io_out_bits_centeroidIndex = T237;
  assign T237 = outputReg_0_centeroidIndex & T238;
  assign T238 = {5'h10/* 16*/{T22}};
  assign io_out_bits_centeroidsFinished = T240;
  assign T240 = outputReg_0_centeroidsFinished & T22;
  assign io_out_bits_point_y = T242;
  assign T242 = outputReg_0_point_y & T243;
  assign T243 = {7'h40/* 64*/{T22}};
  assign T244 = T4 ? T245 : outputReg_0_point_y;
  assign T245 = T246[7'h7f/* 127*/:7'h40/* 64*/];
  assign T246 = 192'h0/* 0*/ | T247;
  assign T247 = pMemOut_0_rData & T248;
  assign T248 = {8'hc0/* 192*/{T5}};
  assign T249 = T250 || T4;
  assign T250 = T180 || T251;
  assign T251 = T154 && T5;
  assign T252 = T338 ? T253 : pMemOut_0_rData;
  assign T253 = partialAccumulatorMemPortReplyValue[8'hbf/* 191*/:1'h0/* 0*/];
  assign partialAccumulatorMemPortReplyValue = T335 ? T334 : T254;
  assign T254 = {T255};
  assign T255 = partialAccumulatorMemPortReplyStorage_0_rData & T256;
  assign T256 = {8'hc0/* 192*/{T5}};
  assign T257 = partialAccumulatorMemPort_rep_valid && T258;
  assign T258 = T259;
  assign T259 = T260[1'h0/* 0*/:1'h0/* 0*/];
  assign T260 = 1'h1/* 1*/ << partialAccumulatorMemPort_rep_tag;
  assign T261 = T257 ? partialAccumulatorMemPort_rep_bits_rData : partialAccumulatorMemPortReplyStorage_0_rData;
  assign partialAccumulatorMemPort_rep_bits_rData = mainOff_partialAccumulatorMem_rep_bits_rData;
  assign mainOff_partialAccumulatorMem_req_bits_wData = partialAccumulatorMemPort_req_bits_wData;
  assign partialAccumulatorMemPort_req_bits_wData = T262;
  assign T262 = T263[8'hc0/* 192*/:1'h1/* 1*/];
  assign T263 = T328 ? T326 : T264;
  assign T264 = {T325, T324, T323, T265};
  assign T265 = T266[1'h0/* 0*/];
  assign T266 = T319 ? T281 : T267;
  assign T267 = {T280, T279, T278, T268};
  assign T268 = T269[1'h0/* 0*/];
  assign T269 = T274 ? T271 : T270;
  assign T270 = {194'h0/* 0*/, 32'h0/* 0*/};
  assign T271 = {pMemIn3_addr, pMemIn3_rw, pMemIn3_wData, pMemIn3_initialize};
  assign pMemIn3_rw = 1'h0/* 0*/;
  assign pMemIn3_addr = T272;
  assign T272 = centeroidIndex_0 & T273;
  assign T273 = {6'h20/* 32*/{T22}};
  assign T274 = T277 && T275;
  assign T275 = T20 == T276;
  assign T276 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign T277 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T278 = T269[8'hc0/* 192*/:1'h1/* 1*/];
  assign T279 = T269[8'hc1/* 193*/];
  assign T280 = T269[8'he1/* 225*/:8'hc2/* 194*/];
  assign T281 = {pMemIn2_addr, pMemIn2_rw, pMemIn2_wData, pMemIn2_initialize};
  assign pMemIn2_wData = T282;
  assign T282 = 192'h0/* 0*/ | T283;
  assign T283 = {T310, T304, T284};
  assign T284 = memData_0_z & T285;
  assign T285 = {7'h40/* 64*/{T22}};
  assign T286 = T174 || T162;
  assign T287 = T162 ? addOut3_out : T288;
  assign T288 = T174 ? T289 : memData_0_z;
  assign T289 = T290[6'h3f/* 63*/:1'h0/* 0*/];
  assign T290 = 192'h0/* 0*/ | T247;
  assign addOut3_out = T291;
  assign T291 = addPortReplyValue[6'h3f/* 63*/:1'h0/* 0*/];
  assign addPortReplyValue = T301 ? T300 : T292;
  assign T292 = {T293};
  assign T293 = addPortReplyStorage_0_out & T294;
  assign T294 = {7'h40/* 64*/{T5}};
  assign T295 = addPort_rep_valid && T296;
  assign T296 = T297;
  assign T297 = T298[1'h0/* 0*/:1'h0/* 0*/];
  assign T298 = 1'h1/* 1*/ << addPort_rep_tag;
  assign T299 = T295 ? addPort_rep_bits_out : addPortReplyStorage_0_out;
  assign addPort_rep_bits_out = mainOff_add_rep_bits_out;
  assign T300 = {addPort_rep_bits_out};
  assign T301 = addPort_rep_valid && T302;
  assign T302 = T303 == addPort_rep_tag;
  assign T303 = {9'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T304 = memData_0_y & T305;
  assign T305 = {7'h40/* 64*/{T22}};
  assign T306 = T174 || T168;
  assign T307 = T168 ? addOut2_out : T308;
  assign T308 = T174 ? T309 : memData_0_y;
  assign T309 = T290[7'h7f/* 127*/:7'h40/* 64*/];
  assign addOut2_out = T291;
  assign T310 = memData_0_x & T311;
  assign T311 = {7'h40/* 64*/{T22}};
  assign T312 = T174 || T174;
  assign T313 = T174 ? addOut1_out : T314;
  assign T314 = T174 ? T315 : memData_0_x;
  assign T315 = T290[8'hbf/* 191*/:8'h80/* 128*/];
  assign addOut1_out = T291;
  assign pMemIn2_rw = 1'h1/* 1*/;
  assign pMemIn2_addr = T316;
  assign T316 = {16'h0/* 0*/, T317};
  assign T317 = inputReg_0_centeroidIndex & T318;
  assign T318 = {5'h10/* 16*/{T22}};
  assign T319 = T322 && T320;
  assign T320 = T20 == T321;
  assign T321 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign T322 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign T323 = T266[8'hc0/* 192*/:1'h1/* 1*/];
  assign T324 = T266[8'hc1/* 193*/];
  assign T325 = T266[8'he1/* 225*/:8'hc2/* 194*/];
  assign T326 = {pMemIn1_addr, pMemIn1_rw, pMemIn1_wData, pMemIn1_initialize};
  assign pMemIn1_rw = 1'h0/* 0*/;
  assign pMemIn1_addr = T327;
  assign T327 = {16'h0/* 0*/, T317};
  assign T328 = T331 && T329;
  assign T329 = T20 == T330;
  assign T330 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign T331 = rThreadEncoder_io_chosen != 1'h1/* 1*/;
  assign mainOff_partialAccumulatorMem_req_bits_addr = partialAccumulatorMemPort_req_bits_addr;
  assign partialAccumulatorMemPort_req_bits_addr = T332;
  assign T332 = T263[8'he1/* 225*/:8'hc2/* 194*/];
  assign mainOff_partialAccumulatorMem_req_bits_rw = partialAccumulatorMemPort_req_bits_rw;
  assign partialAccumulatorMemPort_req_bits_rw = T333;
  assign T333 = T263[8'hc1/* 193*/];
  assign T334 = {partialAccumulatorMemPort_rep_bits_rData};
  assign T335 = partialAccumulatorMemPort_rep_valid && T336;
  assign T336 = T337 == partialAccumulatorMemPort_rep_tag;
  assign T337 = {9'h0/* 0*/, vThreadEncoder_io_chosen};
  assign T338 = T339 || T4;
  assign T339 = T180 || T251;
  assign io_out_bits_point_z = T340;
  assign T340 = outputReg_0_point_z & T341;
  assign T341 = {7'h40/* 64*/{T22}};
  assign T342 = T4 ? T343 : outputReg_0_point_z;
  assign T343 = T246[6'h3f/* 63*/:1'h0/* 0*/];
  assign io_out_bits_point_x = T344;
  assign T344 = outputReg_0_point_x & T345;
  assign T345 = {7'h40/* 64*/{T22}};
  assign T346 = T4 ? T347 : outputReg_0_point_x;
  assign T347 = T246[8'hbf/* 191*/:8'h80/* 128*/];
  RREncode_63 rThreadEncoder(
       .io_valid_0( T25 ),
       .io_chosen( rThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_64 vThreadEncoder(
       .io_valid_0( T8 ),
       .io_chosen( vThreadEncoder_io_chosen ),
       .io_ready(  ));
  RREncode_65 sThreadEncoder(
       .io_valid_0( T1 ),
       .io_chosen( sThreadEncoder_io_chosen ),
       .io_ready(  ));

  always @(posedge clk) begin
    if(reset) begin
      State_0 <= 8'h0/* 0*/;
    end else if(T3) begin
      State_0 <= T191;
    end
    addPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T12;
    subStateTh_0 <= reset ? 1'h0/* 0*/ : T26;
    addPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T40;
    add_ready_received <= reset ? 1'h0/* 0*/ : T44;
    partialAccumulatorMem_valid_received_0 <= reset ? 1'h0/* 0*/ : T68;
    partialAccumulatorMemPortHadReadyRequest <= reset ? 1'h0/* 0*/ : T79;
    partialAccumulatorMem_ready_received <= reset ? 1'h0/* 0*/ : T83;
    add_valid_received_0 <= reset ? 1'h0/* 0*/ : T99;
    partialAccumulatorMemPortHadValidRequest_0 <= reset ? 1'h0/* 0*/ : T120;
    if(T147) begin
      inputReg_0_centeroidIndex <= T153;
    end
    if(reset) begin
      EmitReturnState_0 <= 8'h0/* 0*/;
    end else if(T203) begin
      EmitReturnState_0 <= T220;
    end
    if(reset) begin
      centeroidIndex_0 <= 32'h0/* 0*/;
    end else if(T210) begin
      centeroidIndex_0 <= T215;
    end
    if(T147) begin
      inputTag_0 <= T231;
    end
    outputReg_0_pointsFinished <= T236;
    outputReg_0_centeroidIndex <= T239;
    outputReg_0_centeroidsFinished <= T241;
    if(T4) begin
      outputReg_0_point_y <= T244;
    end
    if(T249) begin
      pMemOut_0_rData <= T252;
    end
    if(T257) begin
      partialAccumulatorMemPortReplyStorage_0_rData <= T261;
    end
    if(T286) begin
      memData_0_z <= T287;
    end
    if(T295) begin
      addPortReplyStorage_0_out <= T299;
    end
    if(T306) begin
      memData_0_y <= T307;
    end
    if(T312) begin
      memData_0_x <= T313;
    end
    if(T4) begin
      outputReg_0_point_z <= T342;
    end
    if(T4) begin
      outputReg_0_point_x <= T346;
    end
  end
endmodule

module rawSpMem_20(input clk, input reset,
    input [9:0] io_addr,
    input  io_rw,
    input [191:0] io_wData,
    output[191:0] io_rData);

  wire[191:0] T0;
  reg [191:0] ram [999:0];
  wire[191:0] T1;
  wire[191:0] T2;
  wire T3;
  wire[191:0] T4;
  wire[9:0] T5;
  reg[191:0] rAddrReg;
  wire[9:0] T6;

  assign io_rData = T0;
  assign T0 = ram[T6];
  assign T2 = io_wData;
  assign T3 = io_rw == 1'h1/* 1*/;
  assign T5 = rAddrReg[4'h9/* 9*/:1'h0/* 0*/];
  assign T6 = rAddrReg[4'h9/* 9*/:1'h0/* 0*/];

  always @(posedge clk) begin
    if (T3)
      ram[io_addr] <= T2;
    rAddrReg <= io_addr;
  end
endmodule

module spMemComponent_20(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [9:0] io_in_bits_addr,
    input  io_in_bits_rw,
    input [191:0] io_in_bits_wData,
    input  io_in_bits_initialize,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[191:0] io_out_bits_rData,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  reg[9:0] tagReg;
  reg[0:0] hasReqReg;
  wire[191:0] rspm_io_rData;

  assign io_out_tag = tagReg;
  assign io_out_valid = hasReqReg;
  assign io_in_ready = io_out_ready;
  assign io_out_bits_rData = rspm_io_rData;
  rawSpMem_20 rspm(.clk(clk), .reset(reset),
       .io_addr( io_in_bits_addr ),
       .io_rw( io_in_bits_rw ),
       .io_wData( io_in_bits_wData ),
       .io_rData( rspm_io_rData ));

  always @(posedge clk) begin
    tagReg <= io_in_tag;
    hasReqReg <= reset ? 1'h0/* 0*/ : io_in_valid;
  end
endmodule

module gOffloadedComponent_130(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType,
    input  mainOff_add_req_ready,
    output mainOff_add_req_valid,
    output[63:0] mainOff_add_req_bits_in1,
    output[63:0] mainOff_add_req_bits_in2,
    output[9:0] mainOff_add_req_tag,
    output mainOff_add_rep_ready,
    input  mainOff_add_rep_valid,
    input [63:0] mainOff_add_rep_bits_out,
    input [9:0] mainOff_add_rep_tag);

  wire mainComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_partialAccumulatorMem_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_partialAccumulatorMem_req_valid;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_partialAccumulatorMem_rep_ready;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;
  wire mainComp_io_out_bits_pointsFinished;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire mainComp_io_out_bits_centeroidsFinished;
  wire[63:0] mainComp_io_out_bits_point_y;
  wire[191:0] offComp_io_out_bits_rData;
  wire[191:0] mainComp_mainOff_partialAccumulatorMem_req_bits_wData;
  wire[9:0] T0;
  wire[31:0] mainComp_mainOff_partialAccumulatorMem_req_bits_addr;
  wire mainComp_mainOff_partialAccumulatorMem_req_bits_rw;
  wire[63:0] mainComp_io_out_bits_point_z;
  wire[63:0] mainComp_io_out_bits_point_x;

  assign io_in_ready = mainComp_io_in_ready;
  assign mainOff_add_rep_ready = mainComp_mainOff_add_rep_ready;
  assign mainOff_add_req_tag = mainComp_mainOff_add_req_tag;
  assign mainOff_add_req_valid = mainComp_mainOff_add_req_valid;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_pointsFinished = mainComp_io_out_bits_pointsFinished;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_bits_centeroidsFinished = mainComp_io_out_bits_centeroidsFinished;
  assign io_out_bits_point_y = mainComp_io_out_bits_point_y;
  assign T0 = mainComp_mainOff_partialAccumulatorMem_req_bits_addr[4'h9/* 9*/:1'h0/* 0*/];
  assign io_out_bits_point_z = mainComp_io_out_bits_point_z;
  assign io_out_bits_point_x = mainComp_io_out_bits_point_x;
  KReduce mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished(  ),
       .io_in_bits_pointsFinished(  ),
       .io_in_bits_centeroidIndex( io_in_bits_centeroidIndex ),
       .io_in_bits_point_x(  ),
       .io_in_bits_point_y(  ),
       .io_in_bits_point_z(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished( mainComp_io_out_bits_centeroidsFinished ),
       .io_out_bits_pointsFinished( mainComp_io_out_bits_pointsFinished ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x( mainComp_io_out_bits_point_x ),
       .io_out_bits_point_y( mainComp_io_out_bits_point_y ),
       .io_out_bits_point_z( mainComp_io_out_bits_point_z ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_partialAccumulatorMem_req_ready( offComp_io_in_ready ),
       .mainOff_partialAccumulatorMem_req_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .mainOff_partialAccumulatorMem_req_bits_addr( mainComp_mainOff_partialAccumulatorMem_req_bits_addr ),
       .mainOff_partialAccumulatorMem_req_bits_rw( mainComp_mainOff_partialAccumulatorMem_req_bits_rw ),
       .mainOff_partialAccumulatorMem_req_bits_wData( mainComp_mainOff_partialAccumulatorMem_req_bits_wData ),
       .mainOff_partialAccumulatorMem_req_bits_initialize(  ),
       .mainOff_partialAccumulatorMem_req_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .mainOff_partialAccumulatorMem_rep_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .mainOff_partialAccumulatorMem_rep_valid( offComp_io_out_valid ),
       .mainOff_partialAccumulatorMem_rep_bits_rData( offComp_io_out_bits_rData ),
       .mainOff_partialAccumulatorMem_rep_tag( offComp_io_out_tag ),
       .mainOff_add_req_ready( mainOff_add_req_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1(  ),
       .mainOff_add_req_bits_in2(  ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( mainOff_add_rep_valid ),
       .mainOff_add_rep_bits_out( mainOff_add_rep_bits_out ),
       .mainOff_add_rep_tag( mainOff_add_rep_tag ));
  spMemComponent_20 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_partialAccumulatorMem_req_valid ),
       .io_in_bits_addr( T0 ),
       .io_in_bits_rw( mainComp_mainOff_partialAccumulatorMem_req_bits_rw ),
       .io_in_bits_wData( mainComp_mainOff_partialAccumulatorMem_req_bits_wData ),
       .io_in_bits_initialize(  ),
       .io_in_tag( mainComp_mainOff_partialAccumulatorMem_req_tag ),
       .io_out_ready( mainComp_mainOff_partialAccumulatorMem_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits_rData( offComp_io_out_bits_rData ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gPipe_100(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [31:0] io_in_bits,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire[9:0] T0;
  reg[4:0] tags_3;
  reg[4:0] tags_2;
  reg[4:0] tags_1;
  reg[4:0] tags_0;
  reg[0:0] valids_3;
  reg[0:0] valids_2;
  reg[0:0] valids_1;
  reg[0:0] valids_0;

  assign io_in_ready = io_out_ready;
  assign io_out_tag = T0;
  assign T0 = {5'h0/* 0*/, tags_3};
  assign io_out_valid = valids_3;

  always @(posedge clk) begin
    if(io_out_ready) begin
      tags_3 <= tags_2;
    end
    if(io_out_ready) begin
      tags_2 <= tags_1;
    end
    if(io_out_ready) begin
      tags_1 <= tags_0;
    end
    if(io_out_ready) begin
      tags_0 <= io_in_tag;
    end
    if(reset) begin
      valids_3 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_3 <= valids_2;
    end
    if(reset) begin
      valids_2 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_2 <= valids_1;
    end
    if(reset) begin
      valids_1 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_1 <= valids_0;
    end
    if(reset) begin
      valids_0 <= 1'h0/* 0*/;
    end else if(io_out_ready) begin
      valids_0 <= io_in_valid;
    end
  end
endmodule

module FUSynWrapper_100(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [63:0] io_in_bits_in1,
    input [63:0] io_in_bits_in2,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output[63:0] io_out_bits,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire tagPipe_io_in_ready;
  wire[9:0] tagPipe_io_out_tag;
  wire T0;
  wire tagPipe_io_out_valid;
  wire bb_io_rdy;

  assign io_in_ready = tagPipe_io_in_ready;
  assign io_out_tag = tagPipe_io_out_tag;
  assign io_out_valid = T0;
  assign T0 = bb_io_rdy && tagPipe_io_out_valid;
  assign T1 = 1'h1/* 1*/;
  gPipe_100 tagPipe(.clk(clk), .reset(reset),
       .io_in_ready( tagPipe_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits(  ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( tagPipe_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( tagPipe_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  types_float_double_grp_fu_86_ACMP_dadd_2_io bb(
       .io_a( io_in_bits_in1 ),
       .io_b( io_in_bits_in2 ),
       .io_result(  ),
       .io_ce( T1 ),
       .io_rdy( bb_io_rdy ));
endmodule

module gOffloadedComponent_131(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire mainComp_io_in_ready;
  wire offComp_io_in_ready;
  wire mainComp_mainOff_add_rep_ready;
  wire[9:0] offComp_io_out_tag;
  wire[9:0] mainComp_mainOff_add_req_tag;
  wire offComp_io_out_valid;
  wire mainComp_mainOff_add_req_valid;
  wire[9:0] mainComp_io_out_tag;
  wire mainComp_io_out_valid;
  wire mainComp_io_out_bits_pointsFinished;
  wire[15:0] mainComp_io_out_bits_centeroidIndex;
  wire mainComp_io_out_bits_centeroidsFinished;
  wire[63:0] mainComp_io_out_bits_point_y;
  wire[63:0] mainComp_io_out_bits_point_z;
  wire[63:0] mainComp_io_out_bits_point_x;
  wire[63:0] mainComp_mainOff_add_req_bits_in1;
  wire[63:0] mainComp_mainOff_add_req_bits_in2;

  assign io_in_ready = mainComp_io_in_ready;
  assign io_out_tag = mainComp_io_out_tag;
  assign io_out_valid = mainComp_io_out_valid;
  assign io_out_bits_pointsFinished = mainComp_io_out_bits_pointsFinished;
  assign io_out_bits_centeroidIndex = mainComp_io_out_bits_centeroidIndex;
  assign io_out_bits_centeroidsFinished = mainComp_io_out_bits_centeroidsFinished;
  assign io_out_bits_point_y = mainComp_io_out_bits_point_y;
  assign io_out_bits_point_z = mainComp_io_out_bits_point_z;
  assign io_out_bits_point_x = mainComp_io_out_bits_point_x;
  gOffloadedComponent_130 mainComp(.clk(clk), .reset(reset),
       .io_in_ready( mainComp_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished(  ),
       .io_in_bits_pointsFinished(  ),
       .io_in_bits_centeroidIndex( io_in_bits_centeroidIndex ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( mainComp_io_out_valid ),
       .io_out_bits_centeroidsFinished( mainComp_io_out_bits_centeroidsFinished ),
       .io_out_bits_pointsFinished( mainComp_io_out_bits_pointsFinished ),
       .io_out_bits_centeroidIndex( mainComp_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x( mainComp_io_out_bits_point_x ),
       .io_out_bits_point_y( mainComp_io_out_bits_point_y ),
       .io_out_bits_point_z( mainComp_io_out_bits_point_z ),
       .io_out_tag( mainComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ),
       .mainOff_add_req_ready( offComp_io_in_ready ),
       .mainOff_add_req_valid( mainComp_mainOff_add_req_valid ),
       .mainOff_add_req_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .mainOff_add_req_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .mainOff_add_req_tag( mainComp_mainOff_add_req_tag ),
       .mainOff_add_rep_ready( mainComp_mainOff_add_rep_ready ),
       .mainOff_add_rep_valid( offComp_io_out_valid ),
       .mainOff_add_rep_bits_out(  ),
       .mainOff_add_rep_tag( offComp_io_out_tag ));
  FUSynWrapper_100 offComp(.clk(clk), .reset(reset),
       .io_in_ready( offComp_io_in_ready ),
       .io_in_valid( mainComp_mainOff_add_req_valid ),
       .io_in_bits_in1( mainComp_mainOff_add_req_bits_in1 ),
       .io_in_bits_in2( mainComp_mainOff_add_req_bits_in2 ),
       .io_in_tag( mainComp_mainOff_add_req_tag ),
       .io_out_ready( mainComp_mainOff_add_rep_ready ),
       .io_out_valid( offComp_io_out_valid ),
       .io_out_bits(  ),
       .io_out_tag( offComp_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module gChainedComponent_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire source_io_in_ready;
  wire sink_io_in_ready;
  wire source_io_out_valid;
  wire[15:0] source_io_out_bits_centeroidIndex;
  wire[9:0] sink_io_out_tag;
  wire[9:0] source_io_out_tag;
  wire sink_io_out_valid;
  wire sink_io_out_bits_pointsFinished;
  wire[15:0] sink_io_out_bits_centeroidIndex;
  wire sink_io_out_bits_centeroidsFinished;
  wire[63:0] sink_io_out_bits_point_y;
  wire[63:0] sink_io_out_bits_point_z;
  wire[63:0] sink_io_out_bits_point_x;
  wire[63:0] source_io_out_bits_point_z;
  wire[63:0] source_io_out_bits_point_y;
  wire[63:0] source_io_out_bits_point_x;

  assign io_in_ready = source_io_in_ready;
  assign io_out_tag = sink_io_out_tag;
  assign io_out_valid = sink_io_out_valid;
  assign io_out_bits_pointsFinished = sink_io_out_bits_pointsFinished;
  assign io_out_bits_centeroidIndex = sink_io_out_bits_centeroidIndex;
  assign io_out_bits_centeroidsFinished = sink_io_out_bits_centeroidsFinished;
  assign io_out_bits_point_y = sink_io_out_bits_point_y;
  assign io_out_bits_point_z = sink_io_out_bits_point_z;
  assign io_out_bits_point_x = sink_io_out_bits_point_x;
  gChainedComponent source(.clk(clk), .reset(reset),
       .io_in_ready( source_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( sink_io_in_ready ),
       .io_out_valid( source_io_out_valid ),
       .io_out_bits_centeroidsFinished(  ),
       .io_out_bits_pointsFinished(  ),
       .io_out_bits_centeroidIndex( source_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x( source_io_out_bits_point_x ),
       .io_out_bits_point_y( source_io_out_bits_point_y ),
       .io_out_bits_point_z( source_io_out_bits_point_z ),
       .io_out_tag( source_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
  gOffloadedComponent_131 sink(.clk(clk), .reset(reset),
       .io_in_ready( sink_io_in_ready ),
       .io_in_valid( source_io_out_valid ),
       .io_in_bits_centeroidsFinished(  ),
       .io_in_bits_pointsFinished(  ),
       .io_in_bits_centeroidIndex( source_io_out_bits_centeroidIndex ),
       .io_in_bits_point_x( source_io_out_bits_point_x ),
       .io_in_bits_point_y( source_io_out_bits_point_y ),
       .io_in_bits_point_z( source_io_out_bits_point_z ),
       .io_in_tag( source_io_out_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( sink_io_out_valid ),
       .io_out_bits_centeroidsFinished( sink_io_out_bits_centeroidsFinished ),
       .io_out_bits_pointsFinished( sink_io_out_bits_pointsFinished ),
       .io_out_bits_centeroidIndex( sink_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x( sink_io_out_bits_point_x ),
       .io_out_bits_point_y( sink_io_out_bits_point_y ),
       .io_out_bits_point_z( sink_io_out_bits_point_z ),
       .io_out_tag( sink_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

module Top(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input  io_in_bits_centeroidsFinished,
    input  io_in_bits_pointsFinished,
    input [15:0] io_in_bits_centeroidIndex,
    input [63:0] io_in_bits_point_x,
    input [63:0] io_in_bits_point_y,
    input [63:0] io_in_bits_point_z,
    input [9:0] io_in_tag,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_centeroidsFinished,
    output io_out_bits_pointsFinished,
    output[15:0] io_out_bits_centeroidIndex,
    output[63:0] io_out_bits_point_x,
    output[63:0] io_out_bits_point_y,
    output[63:0] io_out_bits_point_z,
    output[9:0] io_out_tag,
    input  io_pcIn_valid,
    input  io_pcIn_bits_request,
    input [15:0] io_pcIn_bits_moduleId,
    input [7:0] io_pcIn_bits_portId,
    input [19:0] io_pcIn_bits_pcValue,
    input [3:0] io_pcIn_bits_pcType,
    output io_pcOut_valid,
    output io_pcOut_bits_request,
    output[15:0] io_pcOut_bits_moduleId,
    output[7:0] io_pcOut_bits_portId,
    output[19:0] io_pcOut_bits_pcValue,
    output[3:0] io_pcOut_bits_pcType);

  wire generatedTop_io_in_ready;
  wire[9:0] generatedTop_io_out_tag;
  wire generatedTop_io_out_valid;
  wire generatedTop_io_out_bits_pointsFinished;
  wire[15:0] generatedTop_io_out_bits_centeroidIndex;
  wire generatedTop_io_out_bits_centeroidsFinished;
  wire[63:0] generatedTop_io_out_bits_point_y;
  wire[63:0] generatedTop_io_out_bits_point_z;
  wire[63:0] generatedTop_io_out_bits_point_x;

  assign io_in_ready = generatedTop_io_in_ready;
  assign io_out_tag = generatedTop_io_out_tag;
  assign io_out_valid = generatedTop_io_out_valid;
  assign io_out_bits_pointsFinished = generatedTop_io_out_bits_pointsFinished;
  assign io_out_bits_centeroidIndex = generatedTop_io_out_bits_centeroidIndex;
  assign io_out_bits_centeroidsFinished = generatedTop_io_out_bits_centeroidsFinished;
  assign io_out_bits_point_y = generatedTop_io_out_bits_point_y;
  assign io_out_bits_point_z = generatedTop_io_out_bits_point_z;
  assign io_out_bits_point_x = generatedTop_io_out_bits_point_x;
  gChainedComponent_1 generatedTop(.clk(clk), .reset(reset),
       .io_in_ready( generatedTop_io_in_ready ),
       .io_in_valid( io_in_valid ),
       .io_in_bits_centeroidsFinished( io_in_bits_centeroidsFinished ),
       .io_in_bits_pointsFinished( io_in_bits_pointsFinished ),
       .io_in_bits_centeroidIndex(  ),
       .io_in_bits_point_x( io_in_bits_point_x ),
       .io_in_bits_point_y( io_in_bits_point_y ),
       .io_in_bits_point_z( io_in_bits_point_z ),
       .io_in_tag( io_in_tag ),
       .io_out_ready( io_out_ready ),
       .io_out_valid( generatedTop_io_out_valid ),
       .io_out_bits_centeroidsFinished( generatedTop_io_out_bits_centeroidsFinished ),
       .io_out_bits_pointsFinished( generatedTop_io_out_bits_pointsFinished ),
       .io_out_bits_centeroidIndex( generatedTop_io_out_bits_centeroidIndex ),
       .io_out_bits_point_x( generatedTop_io_out_bits_point_x ),
       .io_out_bits_point_y( generatedTop_io_out_bits_point_y ),
       .io_out_bits_point_z( generatedTop_io_out_bits_point_z ),
       .io_out_tag( generatedTop_io_out_tag ),
       .io_pcIn_valid(  ),
       .io_pcIn_bits_request(  ),
       .io_pcIn_bits_moduleId(  ),
       .io_pcIn_bits_portId(  ),
       .io_pcIn_bits_pcValue(  ),
       .io_pcIn_bits_pcType(  ),
       .io_pcOut_valid(  ),
       .io_pcOut_bits_request(  ),
       .io_pcOut_bits_moduleId(  ),
       .io_pcOut_bits_portId(  ),
       .io_pcOut_bits_pcValue(  ),
       .io_pcOut_bits_pcType(  ));
endmodule

